----------------------------------------------------------------------------------
-- Company: DHBW
-- Engineer: 
-- 
-- Create Date: 05/23/2021 11:12:41 AM
-- Design Name: 
-- Module Name: 
-- Project Name: EDRICO
-- Target Devices: Arty Z7
-- Tool Versions: 
-- Description: 
--  this package contains stimuli and verification dat for the 
--  .vhd testbench.
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


----------------------------------------------------------------------------------
--PACKAGE
----------------------------------------------------------------------------------
package sim_RV32I_RF_UV_1_pkg is
----------------------------------------------------------------------------------
--types
----------------------------------------------------------------------------------
--control_stim(14 downto 10) = register_write, control_stim(9 downto 5) = register_read_A, control_stim(4 downto 0) = register_read_B
type control_stim is array(natural range <>) of std_logic_vector(14 downto 0);
type data_stim  is array(natural range <>) of std_logic_vector(31 downto 0);

--result_vect(63 downto 32)=data_bus_A, result_vect(31 downto 0)=data_bus_B
type result_vect is array(natural range <>) of std_logic_vector(63 downto 0);

----------------------------------------------------------------------------------
--constants
----------------------------------------------------------------------------------
constant results : result_vect(63 downto 0) := 
    (
    0 => x"00000000" & x"00000000",
    1 => x"00000000" & x"00000000",
    2 => x"00000000" & x"00000000",
    3 => x"00000000" & x"00000000",
    4 => x"00000000" & x"00000000",
    5 => x"00000000" & x"00000000",
    6 => x"00000000" & x"00000000",
    7 => x"00000000" & x"00000000",
    8 => x"00000000" & x"00000000",
    9 => x"00000000" & x"00000000",
    10 => x"00000000" & x"00000000",
    11 => x"00000000" & x"00000000",
    12 => x"00000000" & x"00000000",
    13 => x"00000000" & x"00000000",
    14 => x"00000000" & x"00000000",
    15 => x"00000000" & x"00000000",
    16 => x"00000000" & x"00000000",
    17 => x"00000000" & x"00000000",
    18 => x"00000000" & x"00000000",
    19 => x"00000000" & x"00000000",
    20 => x"00000000" & x"00000000",
    21 => x"00000000" & x"00000000",
    22 => x"00000000" & x"00000000",
    23 => x"00000000" & x"00000000",
    24 => x"00000000" & x"00000000",
    25 => x"00000000" & x"00000000",
    26 => x"00000000" & x"00000000",
    27 => x"00000000" & x"00000000",
    28 => x"00000000" & x"00000000",
    29 => x"00000000" & x"00000000",
    30 => x"00000000" & x"00000000",
    31 => x"00000000" & x"00000000",
    32 => x"00000000" & x"00000000",
    33 => x"00000000" & x"00000000",
    34 => x"00000000" & x"00000000",
    35 => x"00000000" & x"00000000",
    36 => x"00000000" & x"00000000",
    37 => x"00000000" & x"00000000",
    38 => x"00000000" & x"00000000",
    39 => x"00000000" & x"00000000",
    40 => x"00000000" & x"00000000",
    41 => x"00000000" & x"00000000",
    42 => x"00000000" & x"00000000",
    43 => x"00000000" & x"00000000",
    44 => x"00000000" & x"00000000",
    45 => x"00000000" & x"00000000",
    46 => x"00000000" & x"00000000",
    47 => x"00000000" & x"00000000",
    48 => x"8BB24E81" & x"0BA73685",
    49 => x"561AC6B1" & x"82364453",
    50 => x"C935C31D" & x"A49A175C",
    51 => x"62E362C9" & x"2B4E1AED",
    52 => x"C819103A" & x"81FC3922",
    53 => x"94168423" & x"C5D219AD",
    54 => x"39381A31" & x"9A892F79",
    55 => x"25624819" & x"ACB390FD",
    56 => x"5F6B51BC" & x"3A8AC9F5",
    57 => x"1BA5864D" & x"369D1CBC",
    58 => x"D4FDA2B0" & x"0C88E6CE",
    59 => x"A3462589" & x"36BD1DEA",
    60 => x"3781B0D4" & x"58311589",
    61 => x"D98BC3A6" & x"8D750715",
    62 => x"48A068DF" & x"F8A00A16",
    63 => x"9F38AA66" & x"00000000"
    );


constant stimulus_data : data_stim(63 downto 0) :=
    (
    0 => x"00000000",
    1 => x"00000000",
    2 => x"00000000",
    3 => x"00000000",
    4 => x"00000000",
    5 => x"00000000",
    6 => x"00000000",
    7 => x"00000000",
    8 => x"00000000",
    9 => x"00000000",
    10 => x"00000000",
    11 => x"00000000",
    12 => x"00000000",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"D7E2E696",
    17 => x"8BB24E81",
    18 => x"0BA73685",
    19 => x"561AC6B1",
    20 => x"82364453",
    21 => x"C935C31D",
    22 => x"A49A175C",
    23 => x"62E362C9",
    24 => x"2B4E1AED",
    25 => x"C819103A",
    26 => x"81FC3922",
    27 => x"94168423",
    28 => x"C5D219AD",
    29 => x"39381A31",
    30 => x"9A892F79",
    31 => x"25624819",
    32 => x"ACB390FD",
    33 => x"5F6B51BC",
    34 => x"3A8AC9F5",
    35 => x"1BA5864D",
    36 => x"369D1CBC",
    37 => x"D4FDA2B0",
    38 => x"0C88E6CE",
    39 => x"A3462589",
    40 => x"36BD1DEA",
    41 => x"3781B0D4",
    42 => x"58311589",
    43 => x"D98BC3A6",
    44 => x"8D750715",
    45 => x"48A068DF",
    46 => x"F8A00A16",
    47 => x"9F38AA66",
    48 => x"00000000",
    49 => x"00000000",
    50 => x"00000000",
    51 => x"00000000",
    52 => x"00000000",
    53 => x"00000000",
    54 => x"00000000",
    55 => x"00000000",
    56 => x"00000000",
    57 => x"00000000",
    58 => x"00000000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000"
    );

constant stimulus_control : control_stim(63 downto 0) :=
    (
    --read all registers after reset(16 cycles)
    0 => "00000" & "00001" & "00010",
    1 => "00000" & "00011" & "00100",
    2 => "00000" & "00101" & "00110",
    3 => "00000" & "00111" & "01000",
    4 => "00000" & "01001" & "01010",
    5 => "00000" & "01011" & "01100",
    6 => "00000" & "01101" & "01110",
    7 => "00000" & "01111" & "10000",
    8 => "00000" & "10001" & "10010",
    9 => "00000" & "10011" & "10100",
    10 => "00000" & "10101" & "10110",
    11 => "00000" & "10111" & "11000",
    12 => "00000" & "11001" & "11010",
    13 => "00000" & "11011" & "11100",
    14 => "00000" & "11101" & "11110",
    15 => "00000" & "11111" & "00000",
    --write to all registers(32 cycles)
    16 => "00000" &	"00000" & "00000",
    17 => "00001" &	"00000" & "00000",
    18 => "00010" &	"00000" & "00000",
    19 => "00011" &	"00000" & "00000",
    20 => "00100" &	"00000" & "00000",
    21 => "00101" &	"00000" & "00000",
    22 => "00110" &	"00000" & "00000",
    23 => "00111" &	"00000" & "00000",
    24 => "01000" &	"00000" & "00000",
    25 => "01001" &	"00000" & "00000",
    26 => "01010" &	"00000" & "00000",
    27 => "01011" &	"00000" & "00000",
    28 => "01100" &	"00000" & "00000",
    29 => "01101" &	"00000" & "00000",
    30 => "01110" &	"00000" & "00000",
    31 => "01111" &	"00000" & "00000",
    32 => "10000" &	"00000" & "00000",
    33 => "10001" &	"00000" & "00000",
    34 => "10010" &	"00000" & "00000",
    35 => "10011" &	"00000" & "00000",
    36 => "10100" &	"00000" & "00000",
    37 => "10101" &	"00000" & "00000",
    38 => "10110" &	"00000" & "00000",
    39 => "10111" &	"00000" & "00000",
    40 => "11000" &	"00000" & "00000",
    41 => "11001" &	"00000" & "00000",
    42 => "11010" &	"00000" & "00000",
    43 => "11011" &	"00000" & "00000",
    44 => "11100" &	"00000" & "00000",
    45 => "11101" &	"00000" & "00000",
    46 => "11110" &	"00000" & "00000",
    47 => "11111" &	"00000" & "00000",
    --read all registers (16 cycles)
    48 => "00000" & "00001" & "00010",
    49 => "00000" & "00011" & "00100",
    50 => "00000" & "00101" & "00110",
    51 => "00000" & "00111" & "01000",
    52 => "00000" & "01001" & "01010",
    53 => "00000" & "01011" & "01100",
    54 => "00000" & "01101" & "01110",
    55 => "00000" & "01111" & "10000",
    56 => "00000" & "10001" & "10010",
    57 => "00000" & "10011" & "10100",
    58 => "00000" & "10101" & "10110",
    59 => "00000" & "10111" & "11000",
    60 => "00000" & "11001" & "11010",
    61 => "00000" & "11011" & "11100",
    62 => "00000" & "11101" & "11110",
    63 => "00000" & "11111" & "00000"
    );



end package;















