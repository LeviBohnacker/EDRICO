----------------------------------------------------------------------------------
-- Company: DHBW
-- Engineer: Levi Bohnacker
-- 
-- Create Date: 05/23/2021 11:12:41 AM
-- Design Name: AXI4_lite_master
-- Module Name: sim_AXI4_CU_UV_2_pkg
-- Project Name: EDRICO
-- Target Devices: Arty Z7
-- Tool Versions: 
-- Description: 
--  this package contains stimuli and verification dat  for the 
--  sim_AXI4_CU_UV_2_tb.vhd testbench.
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


----------------------------------------------------------------------------------
--PACKAGE
----------------------------------------------------------------------------------
package sim_AXI4_CU_UV_2_pkg is
----------------------------------------------------------------------------------
--types
----------------------------------------------------------------------------------
type AXI4_out_rec is record
    --read address channel
    M_AXI_ARCACHE : STD_LOGIC_VECTOR (3 downto 0);
    M_AXI_ARPROT : STD_LOGIC_VECTOR (2 downto 0);
    M_AXI_ARVALID : STD_LOGIC;
    --read data channel
    M_AXI_RREADY : STD_LOGIC;
    --write address channel
    M_AXI_AWCACHE : STD_LOGIC_VECTOR (3 downto 0);
    M_AXI_AWPROT : STD_LOGIC_VECTOR (2 downto 0);
    M_AXI_AWVALID : STD_LOGIC;
    --write data channel
    M_AXI_WSTRB : STD_LOGIC_VECTOR (3 downto 0);
    M_AXI_WVALID : STD_LOGIC;
    --write response channel
    M_AXI_BREADY : STD_LOGIC;
end record AXI4_out_rec;

type AXI4_in_rec is record
    --read address channel
    M_AXI_ARREADY : STD_LOGIC;
    --read data channel
    M_AXI_RRESP : STD_LOGIC_VECTOR (1 downto 0);
    M_AXI_RVALID : STD_LOGIC;
    --write address channel
    M_AXI_AWREADY : STD_LOGIC;
    --write data channel
    M_AXI_WREADY : STD_LOGIC;
    --write response channel
    M_AXI_BRESP : STD_LOGIC_VECTOR (1 downto 0);
    M_AXI_BVALID : STD_LOGIC;
end record AXI4_in_rec;

type input_rec is record
    --controll signals
    enable : STD_LOGIC;
    readWrite : STD_LOGIC;
    instruction : STD_LOGIC;
    size : STD_LOGIC_VECTOR(1 downto 0);
    --halt core
    halt_core : STD_LOGIC;
end record input_rec;

type output_rec is record
    --system control
    memOp_finished : STD_LOGIC;
    store_systemData : STD_LOGIC;
    --exception flags
    load_afe_AXI : STD_LOGIC;
    storeAMO_afe_AXI : STD_LOGIC;
    instruction_afe_AXI : STD_LOGIC;
    --register control
    load_address : STD_LOGIC;
    load_data : STD_LOGIC;
end record output_rec;

type output_vec is array(natural range <>) of output_rec;
type input_vec is array(natural range <>) of input_rec;
type AXI4_in_vec is array(natural range <>) of AXI4_in_rec;
type AXI4_out_vec is array(natural range <>) of AXI4_out_rec;

----------------------------------------------------------------------------------
--constants
----------------------------------------------------------------------------------
constant stimulus_input : input_vec(45 downto 0) := (
    0 => (enable => '0',readWrite => '0',instruction => '0',size => "00",halt_core => '0'),
    --write transfer test
    1 => (enable => '1',readWrite => '1',instruction => '0',size => "10",halt_core => '0'),
    2 => (enable => '1',readWrite => '1',instruction => '0',size => "10",halt_core => '0'),
    3 => (enable => '1',readWrite => '1',instruction => '0',size => "10",halt_core => '0'),
    4 => (enable => '0',readWrite => '0',instruction => '0',size => "00",halt_core => '0'),
    --read transfer test
    5 => (enable => '1',readWrite => '0',instruction => '0',size => "10",halt_core => '0'),
    6 => (enable => '1',readWrite => '0',instruction => '0',size => "10",halt_core => '0'),
    7 => (enable => '1',readWrite => '0',instruction => '0',size => "10",halt_core => '0'),
    8 => (enable => '0',readWrite => '0',instruction => '0',size => "00",halt_core => '0'),
    --read instruction test
    9 => (enable => '1',readWrite => '0',instruction => '1',size => "10",halt_core => '0'),
    10 => (enable => '1',readWrite => '0',instruction => '1',size => "10",halt_core => '0'),
    11 => (enable => '1',readWrite => '0',instruction => '1',size => "10",halt_core => '0'),
    12 => (enable => '0',readWrite => '0',instruction => '0',size => "00",halt_core => '0'),
    --write instruction test
    13 => (enable => '1',readWrite => '1',instruction => '1',size => "10",halt_core => '0'),
    14 => (enable => '1',readWrite => '1',instruction => '1',size => "10",halt_core => '0'),
    15 => (enable => '1',readWrite => '1',instruction => '1',size => "10",halt_core => '0'),
    16 => (enable => '0',readWrite => '0',instruction => '0',size => "00",halt_core => '0'),
    --read halfword test
    17 => (enable => '1',readWrite => '0',instruction => '0',size => "01",halt_core => '0'),
    18 => (enable => '1',readWrite => '0',instruction => '0',size => "01",halt_core => '0'),
    19 => (enable => '1',readWrite => '0',instruction => '0',size => "01",halt_core => '0'),
    20 => (enable => '0',readWrite => '0',instruction => '0',size => "00",halt_core => '0'),
    --write byte test
    21 => (enable => '1',readWrite => '1',instruction => '0',size => "00",halt_core => '0'),
    22 => (enable => '1',readWrite => '1',instruction => '0',size => "00",halt_core => '0'),
    23 => (enable => '1',readWrite => '1',instruction => '0',size => "00",halt_core => '0'),
    24 => (enable => '0',readWrite => '0',instruction => '0',size => "00",halt_core => '0'),
    --load_afe test
    25 => (enable => '1',readWrite => '0',instruction => '0',size => "01",halt_core => '0'),
    26 => (enable => '1',readWrite => '0',instruction => '0',size => "01",halt_core => '0'),
    27 => (enable => '1',readWrite => '0',instruction => '0',size => "01",halt_core => '0'),
    28 => (enable => '0',readWrite => '0',instruction => '0',size => "00",halt_core => '0'),
    29 => (enable => '0',readWrite => '0',instruction => '0',size => "00",halt_core => '0'),
    30 => (enable => '0',readWrite => '0',instruction => '0',size => "00",halt_core => '1'),
    31 => (enable => '0',readWrite => '0',instruction => '0',size => "00",halt_core => '0'),
    --storeAMO_afe test
    32 => (enable => '1',readWrite => '1',instruction => '0',size => "10",halt_core => '0'),
    33 => (enable => '1',readWrite => '1',instruction => '0',size => "10",halt_core => '0'),
    34 => (enable => '1',readWrite => '1',instruction => '0',size => "10",halt_core => '0'),
    35 => (enable => '0',readWrite => '0',instruction => '0',size => "00",halt_core => '0'),
    36 => (enable => '0',readWrite => '0',instruction => '0',size => "00",halt_core => '0'),
    37 => (enable => '0',readWrite => '0',instruction => '0',size => "00",halt_core => '1'),
    38 => (enable => '0',readWrite => '0',instruction => '0',size => "00",halt_core => '0'),
    --instruction_afe test
    39 => (enable => '1',readWrite => '0',instruction => '1',size => "01",halt_core => '0'),
    40 => (enable => '1',readWrite => '0',instruction => '1',size => "01",halt_core => '0'),
    41 => (enable => '1',readWrite => '0',instruction => '1',size => "01",halt_core => '0'),
    42 => (enable => '0',readWrite => '0',instruction => '0',size => "00",halt_core => '0'),
    43 => (enable => '0',readWrite => '0',instruction => '0',size => "00",halt_core => '0'),
    44 => (enable => '0',readWrite => '0',instruction => '0',size => "00",halt_core => '1'),
    45 => (enable => '0',readWrite => '0',instruction => '0',size => "00",halt_core => '0')

);

constant stimulus_AXI4_in: AXI4_in_vec(45 downto 0) := (
    0 => (  M_AXI_ARREADY => '0',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '0',
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0'),
    --write transfer test
    1 => (  M_AXI_ARREADY => '0',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '0',
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0'),
    2 => (  M_AXI_ARREADY => '0',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '0',
            M_AXI_AWREADY => '1',
            M_AXI_WREADY => '1',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '1'),
    3 => (  M_AXI_ARREADY => '0',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '0',
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0'),
    4 => (  M_AXI_ARREADY => '0',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '0',
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0'),
    --read transfer test
    5 => (  M_AXI_ARREADY => '0',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '0', 
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0'),
    6 => (  M_AXI_ARREADY => '1',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '1',
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0'),
    7 => (  M_AXI_ARREADY => '0',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '0',
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0'),
    8 => (  M_AXI_ARREADY => '0',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '0',
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0'),
    --read instruction test
    9 => (  M_AXI_ARREADY => '0',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '0', 
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0'),
    10 => (  M_AXI_ARREADY => '1',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '1',
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0'),
    11 => (  M_AXI_ARREADY => '0',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '0',
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0'),
    12 => (  M_AXI_ARREADY => '0',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '0',
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0'),
    --write instruction test
    13 => (  M_AXI_ARREADY => '0',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '0', 
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0'),
    14 => (  M_AXI_ARREADY => '0',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '0',
            M_AXI_AWREADY => '1',
            M_AXI_WREADY => '1',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '1'),
    15 => (  M_AXI_ARREADY => '0',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '0',
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0'),
    16 => (  M_AXI_ARREADY => '0',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '0',
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0'),
    --read halfword
    17 => (  M_AXI_ARREADY => '0',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '0', 
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0'),
    18 => (  M_AXI_ARREADY => '1',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '1',
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0'),
    19 => (  M_AXI_ARREADY => '0',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '0',
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0'),
    20 => (  M_AXI_ARREADY => '0',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '0',
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0'),
    --write byte
    21 => (  M_AXI_ARREADY => '0',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '0', 
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0'),
    22 => (  M_AXI_ARREADY => '0',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '0',
            M_AXI_AWREADY => '1',
            M_AXI_WREADY => '1',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '1'),
    23 => (  M_AXI_ARREADY => '0',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '0',
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0'),
    24 => (  M_AXI_ARREADY => '0',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '0',
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0'),
    --load_afe_test        
    25 => (  M_AXI_ARREADY => '0',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '0', 
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0'),
    26 => (  M_AXI_ARREADY => '1',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '0',
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0'),
    27 => (  M_AXI_ARREADY => '0',
            M_AXI_RRESP => "10",
            M_AXI_RVALID => '1',
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0'),
    28 => (  M_AXI_ARREADY => '0',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '0',
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0'),
    29 => (  M_AXI_ARREADY => '0',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '0',
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0'),
    30 => (  M_AXI_ARREADY => '0',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '0',
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0'),
    31 => (  M_AXI_ARREADY => '0',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '0',
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0'),
    --storeAMO_afe test        
    32 => (  M_AXI_ARREADY => '0',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '0', 
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0'),
    33 => (  M_AXI_ARREADY => '0',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '0',
            M_AXI_AWREADY => '1',
            M_AXI_WREADY => '1',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0'),
    34 => (  M_AXI_ARREADY => '0',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '0',
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "10",
            M_AXI_BVALID => '1'),
    35 => (  M_AXI_ARREADY => '0',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '0',
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0'),
    36 => (  M_AXI_ARREADY => '0',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '0',
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0'),
    37 => (  M_AXI_ARREADY => '0',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '0',
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0'),
    38 => (  M_AXI_ARREADY => '0',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '0',
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0'),
    --instruction_afe test        
    39 => (  M_AXI_ARREADY => '0',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '0', 
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0'),
    40 => (  M_AXI_ARREADY => '1',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '0',
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0'),
    41 => (  M_AXI_ARREADY => '0',
            M_AXI_RRESP => "10",
            M_AXI_RVALID => '1',
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0'),
    42 => (  M_AXI_ARREADY => '0',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '0',
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0'),
    43 => (  M_AXI_ARREADY => '0',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '0',
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0'),
    44 => (  M_AXI_ARREADY => '0',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '0',
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0'),
    45 => (  M_AXI_ARREADY => '0',
            M_AXI_RRESP => "00",
            M_AXI_RVALID => '0',
            M_AXI_AWREADY => '0',
            M_AXI_WREADY => '0',
            M_AXI_BRESP => "00",
            M_AXI_BVALID => '0')
);

constant results_output: output_vec(45 downto 0) := (
    0 => (  memOp_finished => '0',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '0',
            load_data => '0'),
    --write transfer test
    1 => (  memOp_finished => '0',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '1',
            load_data => '1'),
    2 => (  memOp_finished => '0',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '1',
            load_data => '1'),
    3 => (  memOp_finished => '0',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '1',
            load_data => '1'),
    4 => (  memOp_finished => '1',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '0',
            load_data => '0'),
    --read transfer test
    5 => (  memOp_finished => '0',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '1',
            load_data => '0'),
    6 => (  memOp_finished => '0',
            store_systemData => '1',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '1',
            load_data => '0'),
    7 => (  memOp_finished => '0',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '1',
            load_data => '0'),
    8 => (  memOp_finished => '1',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '0',
            load_data => '0'),
    --read instruction test
    9 => (  memOp_finished => '0',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '1',
            load_data => '0'),
    10 => (  memOp_finished => '0',
            store_systemData => '1',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '1',
            load_data => '0'),
    11 => (  memOp_finished => '0',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '1',
            load_data => '0'),
    12 => (  memOp_finished => '1',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '0',
            load_data => '0'),
    --write instruction test
    13 => (  memOp_finished => '0',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '1',
            load_data => '1'),
    14 => (  memOp_finished => '0',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '1',
            load_data => '1'),
    15 => (  memOp_finished => '0',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '1',
            load_data => '1'),
    16 => (  memOp_finished => '1',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '0',
            load_data => '0'),
    --read halfword test
    17 => (  memOp_finished => '0',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '1',
            load_data => '0'),
    18 => (  memOp_finished => '0',
            store_systemData => '1',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '1',
            load_data => '0'),
    19 => (  memOp_finished => '0',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '1',
            load_data => '0'),
    20 => (  memOp_finished => '1',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '0',
            load_data => '0'),
    --write byte test
    21 => (  memOp_finished => '0',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '1',
            load_data => '1'),
    22 => (  memOp_finished => '0',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '1',
            load_data => '1'),
    23 => (  memOp_finished => '0',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '1',
            load_data => '1'),
    24 => (  memOp_finished => '1',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '0',
            load_data => '0'), 
    --load_afe test
    25 => (  memOp_finished => '0',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '1',
            load_data => '0'),
    26 => (  memOp_finished => '0',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '1',
            load_data => '0'),
    27 => (  memOp_finished => '0',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '1',
            load_data => '0'),
    28 => (  memOp_finished => '0',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '0',
            load_data => '0'),
    29 => (  memOp_finished => '0',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '0',
            load_data => '0'),
    30 => (  memOp_finished => '0',
            store_systemData => '0',
            load_afe_AXI => '1',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '0',
            load_data => '0'),
    31 => (  memOp_finished => '0',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '0',
            load_data => '0'), 
    --storeAMO_afe test
    32 => (  memOp_finished => '0',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '1',
            load_data => '1'),
    33 => (  memOp_finished => '0',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '1',
            load_data => '1'),
    34 => (  memOp_finished => '0',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '1',
            load_data => '1'),
    35 => (  memOp_finished => '0',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '0',
            load_data => '0'),
    36 => (  memOp_finished => '0',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '0',
            load_data => '0'),
    37 => (  memOp_finished => '0',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '1',
            instruction_afe_AXI => '0',
            load_address => '0',
            load_data => '0'),
    38 => (  memOp_finished => '0',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '0',
            load_data => '0'), 
    --instruction_afe test
    39 => (  memOp_finished => '0',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '1',
            load_data => '0'),
    40 => (  memOp_finished => '0',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '1',
            load_data => '0'),
    41 => (  memOp_finished => '0',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '1',
            load_data => '0'),
    42 => (  memOp_finished => '0',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '0',
            load_data => '0'),
    43 => (  memOp_finished => '0',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '0',
            load_data => '0'),
    44 => (  memOp_finished => '0',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '1',
            load_address => '0',
            load_data => '0'),
    45 => (  memOp_finished => '0',
            store_systemData => '0',
            load_afe_AXI => '0',
            storeAMO_afe_AXI => '0',
            instruction_afe_AXI => '0',
            load_address => '0',
            load_data => '0')
           
);

constant results_AXI4_out: AXI4_out_vec(45 downto 0) := (
    0 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "000",
            M_AXI_ARVALID => '0',
            M_AXI_RREADY => '0',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "000",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "0001",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '0'),
    --write transfer test
    1 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "000",
            M_AXI_ARVALID => '0',
            M_AXI_RREADY => '0',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "000",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "1111",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '0'),
    2 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "000",
            M_AXI_ARVALID => '0',
            M_AXI_RREADY => '0',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "000",
            M_AXI_AWVALID => '1',
            M_AXI_WSTRB => "1111",
            M_AXI_WVALID => '1',
            M_AXI_BREADY => '1'),
    3 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "000",
            M_AXI_ARVALID => '0',
            M_AXI_RREADY => '0',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "000",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "1111",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '0'),
    4 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "000",
            M_AXI_ARVALID => '0',
            M_AXI_RREADY => '0',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "000",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "0001",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '0'),
    --read transfer test
    5 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "000",
            M_AXI_ARVALID => '0',
            M_AXI_RREADY => '0',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "000",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "1111",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '0'),
    6 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "000",
            M_AXI_ARVALID => '1',
            M_AXI_RREADY => '1',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "000",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "1111",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '0'),
    7 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "000",
            M_AXI_ARVALID => '0',
            M_AXI_RREADY => '0',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "000",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "1111",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '0'),
    8 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "000",
            M_AXI_ARVALID => '0',
            M_AXI_RREADY => '0',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "000",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "0001",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '0'),
    --read instruction test
    9 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "100",
            M_AXI_ARVALID => '0',
            M_AXI_RREADY => '0',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "100",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "1111",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '0'),
    10 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "100",
            M_AXI_ARVALID => '1',
            M_AXI_RREADY => '1',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "100",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "1111",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '0'),
    11 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "100",
            M_AXI_ARVALID => '0',
            M_AXI_RREADY => '0',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "100",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "1111",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '0'),
    12 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "000",
            M_AXI_ARVALID => '0',
            M_AXI_RREADY => '0',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "000",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "0001",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '0'),
    --write instruction test
    13 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "100",
            M_AXI_ARVALID => '0',
            M_AXI_RREADY => '0',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "100",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "1111",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '0'),
    14 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "100",
            M_AXI_ARVALID => '0',
            M_AXI_RREADY => '0',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "100",
            M_AXI_AWVALID => '1',
            M_AXI_WSTRB => "1111",
            M_AXI_WVALID => '1',
            M_AXI_BREADY => '1'),
    15 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "100",
            M_AXI_ARVALID => '0',
            M_AXI_RREADY => '0',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "100",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "1111",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '0'),
    16 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "000",
            M_AXI_ARVALID => '0',
            M_AXI_RREADY => '0',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "000",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "0001",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '0'),
    --read halfword test
    17 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "000",
            M_AXI_ARVALID => '0',
            M_AXI_RREADY => '0',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "000",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "0011",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '0'),
    18 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "000",
            M_AXI_ARVALID => '1',
            M_AXI_RREADY => '1',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "000",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "0011",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '0'),
    19 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "000",
            M_AXI_ARVALID => '0',
            M_AXI_RREADY => '0',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "000",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "0011",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '0'),
    20 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "000",
            M_AXI_ARVALID => '0',
            M_AXI_RREADY => '0',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "000",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "0001",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '0'),
    --write byte test
    21 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "000",
            M_AXI_ARVALID => '0',
            M_AXI_RREADY => '0',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "000",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "0001",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '0'),
    22 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "000",
            M_AXI_ARVALID => '0',
            M_AXI_RREADY => '0',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "000",
            M_AXI_AWVALID => '1',
            M_AXI_WSTRB => "0001",
            M_AXI_WVALID => '1',
            M_AXI_BREADY => '1'),
    23 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "000",
            M_AXI_ARVALID => '0',
            M_AXI_RREADY => '0',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "000",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "0001",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '0'),
    24 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "000",
            M_AXI_ARVALID => '0',
            M_AXI_RREADY => '0',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "000",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "0001",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '0'),
    --loaf_afe test
    25 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "000",
            M_AXI_ARVALID => '0',
            M_AXI_RREADY => '0',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "000",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "0011",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '0'),
    26 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "000",
            M_AXI_ARVALID => '1',
            M_AXI_RREADY => '1',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "000",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "0011",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '0'),
    27 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "000",
            M_AXI_ARVALID => '0',
            M_AXI_RREADY => '1',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "000",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "0011",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '0'),
    28 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "000",
            M_AXI_ARVALID => '0',
            M_AXI_RREADY => '0',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "000",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "0001",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '0'),
    29 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "000",
            M_AXI_ARVALID => '0',
            M_AXI_RREADY => '0',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "000",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "0001",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '0'),
    30 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "000",
            M_AXI_ARVALID => '0',
            M_AXI_RREADY => '0',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "000",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "0001",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '0'),
    31 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "000",
            M_AXI_ARVALID => '0',
            M_AXI_RREADY => '0',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "000",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "0001",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '0'),
    --storeAMO_afe test
    32 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "000",
            M_AXI_ARVALID => '0',
            M_AXI_RREADY => '0',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "000",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "1111",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '0'),
    33 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "000",
            M_AXI_ARVALID => '0',
            M_AXI_RREADY => '0',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "000",
            M_AXI_AWVALID => '1',
            M_AXI_WSTRB => "1111",
            M_AXI_WVALID => '1',
            M_AXI_BREADY => '1'),
    34 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "000",
            M_AXI_ARVALID => '0',
            M_AXI_RREADY => '0',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "000",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "1111",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '1'),
    35 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "000",
            M_AXI_ARVALID => '0',
            M_AXI_RREADY => '0',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "000",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "0001",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '0'),
    36 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "000",
            M_AXI_ARVALID => '0',
            M_AXI_RREADY => '0',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "000",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "0001",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '0'),
    37 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "000",
            M_AXI_ARVALID => '0',
            M_AXI_RREADY => '0',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "000",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "0001",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '0'),
    38 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "000",
            M_AXI_ARVALID => '0',
            M_AXI_RREADY => '0',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "000",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "0001",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '0'),
    --instruction_afe test
    39 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "100",
            M_AXI_ARVALID => '0',
            M_AXI_RREADY => '0',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "100",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "0011",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '0'),
    40 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "100",
            M_AXI_ARVALID => '1',
            M_AXI_RREADY => '1',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "100",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "0011",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '0'),
    41 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "100",
            M_AXI_ARVALID => '0',
            M_AXI_RREADY => '1',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "100",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "0011",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '0'),
    42 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "000",
            M_AXI_ARVALID => '0',
            M_AXI_RREADY => '0',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "000",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "0001",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '0'),
    43 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "000",
            M_AXI_ARVALID => '0',
            M_AXI_RREADY => '0',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "000",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "0001",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '0'),
    44 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "000",
            M_AXI_ARVALID => '0',
            M_AXI_RREADY => '0',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "000",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "0001",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '0'),
    45 => (  M_AXI_ARCACHE => "0011",
            M_AXI_ARPROT => "000",
            M_AXI_ARVALID => '0',
            M_AXI_RREADY => '0',
            M_AXI_AWCACHE => "0011",
            M_AXI_AWPROT => "000",
            M_AXI_AWVALID => '0',
            M_AXI_WSTRB => "0001",
            M_AXI_WVALID => '0',
            M_AXI_BREADY => '0')
);


end package;
