library IEEE
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity testBench is
end entity;

architecture add_test_name of testBench is
--add component

--add pad names
--bsp: 

begin



end architecture;

