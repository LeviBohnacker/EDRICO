----------------------------------------------------------------------------------
-- Company: DHBW
-- Engineer: 
-- 
-- Create Date: 05/23/2021 11:12:41 AM
-- Design Name: 
-- Module Name: 
-- Project Name: EDRICO
-- Target Devices: Arty Z7
-- Tool Versions: 
-- Description: 
--  this package contains stimuli and verification dat for the 
--  .vhd testbench.
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


----------------------------------------------------------------------------------
--PACKAGE
----------------------------------------------------------------------------------
package _UV_x_pkg is
----------------------------------------------------------------------------------
--types
----------------------------------------------------------------------------------

----------------------------------------------------------------------------------
--constants
----------------------------------------------------------------------------------

end package;
