----------------------------------------------------------------------------------
-- Company: DHBW
-- Engineer: Levi Bohnacker
-- 
-- Create Date: 05/23/2021 11:12:41 AM
-- Design Name: RegisterFile
-- Module Name: CSR_controller
-- Project Name: EDRICO
-- Target Devices: Arty Z7
-- Tool Versions: 
-- Description: 
--  this package contains stimuli and verification dat for the 
--  CSR_controller.vhd testbench.
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


----------------------------------------------------------------------------------
--PACKAGE
----------------------------------------------------------------------------------
package sim_CSR_controller_UV_1_pkg is
----------------------------------------------------------------------------------
--types
----------------------------------------------------------------------------------
--input_stimulus(13) = CSR_write, input_stimulus(12) = CSR_read, input_stimulus(11 downto 0) = CSR_address
type input_stim is array(natural range <>) of std_logic_vector(13 downto 0);
--result_vect(39) = illegal_instruction_exception, result_vect(38 downto 33) = CSR_read_sel, result_vect(32 downto 0) = CSR_write_sel
type result_vect is array(natural range <>) of std_logic_vector(39 downto 0);
----------------------------------------------------------------------------------
--constants
-----------------------------------------------ß-----------------------------------
constant stimulus_input : input_stim(255 downto 0) :=
    (
    0 => "1" & "0" &  x"300",
    1 => "1" & "0" &  x"B82",
    2 => "1" & "0" &  x"304",
    3 => "1" & "0" &  x"305",
    4 => "1" & "0" &  x"320",
    5 => "1" & "0" &  x"340",
    6 => "1" & "0" &  x"341",
    7 => "1" & "0" &  x"342",
    8 => "1" & "0" &  x"343",
    9 => "1" & "0" &  x"344",
    10 => "1" & "0" &  x"3A0",
    11 => "1" & "0" &  x"3A1",
    12 => "1" & "0" &  x"3A2",
    13 => "1" & "0" &  x"3A3",
    14 => "1" & "0" &  x"3B0",
    15 => "1" & "0" &  x"3B1",
    16 => "1" & "0" &  x"3B2",
    17 => "1" & "0" &  x"3B3",
    18 => "1" & "0" &  x"3B4",
    19 => "1" & "0" &  x"3B5",
    20 => "1" & "0" &  x"3B6",
    21 => "1" & "0" &  x"3B7",
    22 => "1" & "0" &  x"3B8",
    23 => "1" & "0" &  x"3B9",
    24 => "1" & "0" &  x"3BA",
    25 => "1" & "0" &  x"3BB",
    26 => "1" & "0" &  x"3BC",
    27 => "1" & "0" &  x"3BD",
    28 => "1" & "0" &  x"3BE",
    29 => "1" & "0" &  x"3BF",
    30 => "1" & "0" &  x"B00",
    31 => "1" & "0" &  x"B02",
    32 => "1" & "0" &  x"B80",
    33 => "1" & "0" &  x"301",
    34 => "1" & "0" &  x"323",
    35 => "1" & "0" &  x"324",
    36 => "1" & "0" &  x"325",
    37 => "1" & "0" &  x"326",
    38 => "1" & "0" &  x"327",
    39 => "1" & "0" &  x"328",
    40 => "1" & "0" &  x"329",
    41 => "1" & "0" &  x"32A",
    42 => "1" & "0" &  x"32B",
    43 => "1" & "0" &  x"32C",
    44 => "1" & "0" &  x"32D",
    45 => "1" & "0" &  x"32E",
    46 => "1" & "0" &  x"32F",
    47 => "1" & "0" &  x"330",
    48 => "1" & "0" &  x"331",
    49 => "1" & "0" &  x"332",
    50 => "1" & "0" &  x"333",
    51 => "1" & "0" &  x"334",
    52 => "1" & "0" &  x"335",
    53 => "1" & "0" &  x"336",
    54 => "1" & "0" &  x"337",
    55 => "1" & "0" &  x"338",
    56 => "1" & "0" &  x"339",
    57 => "1" & "0" &  x"33A",
    58 => "1" & "0" &  x"33B",
    59 => "1" & "0" &  x"33C",
    60 => "1" & "0" &  x"33D",
    61 => "1" & "0" &  x"33E",
    62 => "1" & "0" &  x"33F",
    63 => "1" & "0" &  x"B03",
    64 => "1" & "0" &  x"B04",
    65 => "1" & "0" &  x"B05",
    66 => "1" & "0" &  x"B06",
    67 => "1" & "0" &  x"B07",
    68 => "1" & "0" &  x"B08",
    69 => "1" & "0" &  x"B09",
    70 => "1" & "0" &  x"B0A",
    71 => "1" & "0" &  x"B0B",
    72 => "1" & "0" &  x"B0C",
    73 => "1" & "0" &  x"B0D",
    74 => "1" & "0" &  x"B0E",
    75 => "1" & "0" &  x"B0F",
    76 => "1" & "0" &  x"B10",
    77 => "1" & "0" &  x"B11",
    78 => "1" & "0" &  x"B12",
    79 => "1" & "0" &  x"B13",
    80 => "1" & "0" &  x"B14",
    81 => "1" & "0" &  x"B15",
    82 => "1" & "0" &  x"B16",
    83 => "1" & "0" &  x"B17",
    84 => "1" & "0" &  x"B18",
    85 => "1" & "0" &  x"B19",
    86 => "1" & "0" &  x"B1A",
    87 => "1" & "0" &  x"B1B",
    88 => "1" & "0" &  x"B1C",
    89 => "1" & "0" &  x"B1D",
    90 => "1" & "0" &  x"B1E",
    91 => "1" & "0" &  x"B1F",
    92 => "1" & "0" &  x"B83",
    93 => "1" & "0" &  x"B84",
    94 => "1" & "0" &  x"B85",
    95 => "1" & "0" &  x"B86",
    96 => "1" & "0" &  x"B87",
    97 => "1" & "0" &  x"B88",
    98 => "1" & "0" &  x"B89",
    99 => "1" & "0" &  x"B8A",
    100 => "1" & "0" &  x"B8B",
    101 => "1" & "0" &  x"B8C",
    102 => "1" & "0" &  x"B8D",
    103 => "1" & "0" &  x"B8E",
    104 => "1" & "0" &  x"B8F",
    105 => "1" & "0" &  x"B90",
    106 => "1" & "0" &  x"B91",
    107 => "1" & "0" &  x"B92",
    108 => "1" & "0" &  x"B93",
    109 => "1" & "0" &  x"B94",
    110 => "1" & "0" &  x"B95",
    111 => "1" & "0" &  x"B96",
    112 => "1" & "0" &  x"B97",
    113 => "1" & "0" &  x"B98",
    114 => "1" & "0" &  x"B99",
    115 => "1" & "0" &  x"B9A",
    116 => "1" & "0" &  x"B9B",
    117 => "1" & "0" &  x"B9C",
    118 => "1" & "0" &  x"B9D",
    119 => "1" & "0" &  x"B9E",
    120 => "1" & "0" &  x"B9F",
    121 => "1" & "0" &  x"F11",
    122 => "1" & "0" &  x"F12",
    123 => "1" & "0" &  x"F13",
    124 => "1" & "0" &  x"F14",
    125 => "0" & "1" &  x"300",
    126 => "0" & "1" &  x"B82",
    127 => "0" & "1" &  x"304",
    128 => "0" & "1" &  x"305",
    129 => "0" & "1" &  x"320",
    130 => "0" & "1" &  x"340",
    131 => "0" & "1" &  x"341",
    132 => "0" & "1" &  x"342",
    133 => "0" & "1" &  x"343",
    134 => "0" & "1" &  x"344",
    135 => "0" & "1" &  x"3A0",
    136 => "0" & "1" &  x"3A1",
    137 => "0" & "1" &  x"3A2",
    138 => "0" & "1" &  x"3A3",
    139 => "0" & "1" &  x"3B0",
    140 => "0" & "1" &  x"3B1",
    141 => "0" & "1" &  x"3B2",
    142 => "0" & "1" &  x"3B3",
    143 => "0" & "1" &  x"3B4",
    144 => "0" & "1" &  x"3B5",
    145 => "0" & "1" &  x"3B6",
    146 => "0" & "1" &  x"3B7",
    147 => "0" & "1" &  x"3B8",
    148 => "0" & "1" &  x"3B9",
    149 => "0" & "1" &  x"3BA",
    150 => "0" & "1" &  x"3BB",
    151 => "0" & "1" &  x"3BC",
    152 => "0" & "1" &  x"3BD",
    153 => "0" & "1" &  x"3BE",
    154 => "0" & "1" &  x"3BF",
    155 => "0" & "1" &  x"B00",
    156 => "0" & "1" &  x"B02",
    157 => "0" & "1" &  x"B80",
    158 => "0" & "1" &  x"301",
    159 => "0" & "1" &  x"323",
    160 => "0" & "1" &  x"324",
    161 => "0" & "1" &  x"325",
    162 => "0" & "1" &  x"326",
    163 => "0" & "1" &  x"327",
    164 => "0" & "1" &  x"328",
    165 => "0" & "1" &  x"329",
    166 => "0" & "1" &  x"32A",
    167 => "0" & "1" &  x"32B",
    168 => "0" & "1" &  x"32C",
    169 => "0" & "1" &  x"32D",
    170 => "0" & "1" &  x"32E",
    171 => "0" & "1" &  x"32F",
    172 => "0" & "1" &  x"330",
    173 => "0" & "1" &  x"331",
    174 => "0" & "1" &  x"332",
    175 => "0" & "1" &  x"333",
    176 => "0" & "1" &  x"334",
    177 => "0" & "1" &  x"335",
    178 => "0" & "1" &  x"336",
    179 => "0" & "1" &  x"337",
    180 => "0" & "1" &  x"338",
    181 => "0" & "1" &  x"339",
    182 => "0" & "1" &  x"33A",
    183 => "0" & "1" &  x"33B",
    184 => "0" & "1" &  x"33C",
    185 => "0" & "1" &  x"33D",
    186 => "0" & "1" &  x"33E",
    187 => "0" & "1" &  x"33F",
    188 => "0" & "1" &  x"B03",
    189 => "0" & "1" &  x"B04",
    190 => "0" & "1" &  x"B05",
    191 => "0" & "1" &  x"B06",
    192 => "0" & "1" &  x"B07",
    193 => "0" & "1" &  x"B08",
    194 => "0" & "1" &  x"B09",
    195 => "0" & "1" &  x"B0A",
    196 => "0" & "1" &  x"B0B",
    197 => "0" & "1" &  x"B0C",
    198 => "0" & "1" &  x"B0D",
    199 => "0" & "1" &  x"B0E",
    200 => "0" & "1" &  x"B0F",
    201 => "0" & "1" &  x"B10",
    202 => "0" & "1" &  x"B11",
    203 => "0" & "1" &  x"B12",
    204 => "0" & "1" &  x"B13",
    205 => "0" & "1" &  x"B14",
    206 => "0" & "1" &  x"B15",
    207 => "0" & "1" &  x"B16",
    208 => "0" & "1" &  x"B17",
    209 => "0" & "1" &  x"B18",
    210 => "0" & "1" &  x"B19",
    211 => "0" & "1" &  x"B1A",
    212 => "0" & "1" &  x"B1B",
    213 => "0" & "1" &  x"B1C",
    214 => "0" & "1" &  x"B1D",
    215 => "0" & "1" &  x"B1E",
    216 => "0" & "1" &  x"B1F",
    217 => "0" & "1" &  x"B83",
    218 => "0" & "1" &  x"B84",
    219 => "0" & "1" &  x"B85",
    220 => "0" & "1" &  x"B86",
    221 => "0" & "1" &  x"B87",
    222 => "0" & "1" &  x"B88",
    223 => "0" & "1" &  x"B89",
    224 => "0" & "1" &  x"B8A",
    225 => "0" & "1" &  x"B8B",
    226 => "0" & "1" &  x"B8C",
    227 => "0" & "1" &  x"B8D",
    228 => "0" & "1" &  x"B8E",
    229 => "0" & "1" &  x"B8F",
    230 => "0" & "1" &  x"B90",
    231 => "0" & "1" &  x"B91",
    232 => "0" & "1" &  x"B92",
    233 => "0" & "1" &  x"B93",
    234 => "0" & "1" &  x"B94",
    235 => "0" & "1" &  x"B95",
    236 => "0" & "1" &  x"B96",
    237 => "0" & "1" &  x"B97",
    238 => "0" & "1" &  x"B98",
    239 => "0" & "1" &  x"B99",
    240 => "0" & "1" &  x"B9A",
    241 => "0" & "1" &  x"B9B",
    242 => "0" & "1" &  x"B9C",
    243 => "0" & "1" &  x"B9D",
    244 => "0" & "1" &  x"B9E",
    245 => "0" & "1" &  x"B9F",
    246 => "0" & "1" &  x"F11",
    247 => "0" & "1" &  x"F12",
    248 => "0" & "1" &  x"F13",
    249 => "0" & "1" &  x"F14",
    250 => "1" & "1" &  x"FFF",
    251 => "1" & "1" &  x"DEA",
    252 => "1" & "0" &  x"754",
    253 => "0" & "1" &  x"193",
    254 => "0" & "0" &  x"C23",
    255 => "0" & "1" &  x"897" 
    );

constant results : result_vect(255 downto 0) :=
    (
    0 => '0' & "000000" &  '0' & x"00000001",
    1 => '0' & "000000" &  '0' & x"00000002",
    2 => '0' & "000000" &  '0' & x"00000004",
    3 => '0' & "000000" &  '0' & x"00000008",
    4 => '0' & "000000" &  '0' & x"00000010",
    5 => '0' & "000000" &  '0' & x"00000020",
    6 => '0' & "000000" &  '0' & x"00000040",
    7 => '0' & "000000" &  '0' & x"00000080",
    8 => '0' & "000000" &  '0' & x"00000100",
    9 => '0' & "000000" &  '0' & x"00000200",
    10 => '0' & "000000" &  '0' & x"00000400",
    11 => '0' & "000000" &  '0' & x"00000800",
    12 => '0' & "000000" &  '0' & x"00001000",
    13 => '0' & "000000" &  '0' & x"00002000",
    14 => '0' & "000000" &  '0' & x"00004000",
    15 => '0' & "000000" &  '0' & x"00008000",
    16 => '0' & "000000" &  '0' & x"00010000",
    17 => '0' & "000000" &  '0' & x"00020000",
    18 => '0' & "000000" &  '0' & x"00040000",
    19 => '0' & "000000" &  '0' & x"00080000",
    20 => '0' & "000000" &  '0' & x"00100000",
    21 => '0' & "000000" &  '0' & x"00200000",
    22 => '0' & "000000" &  '0' & x"00400000",
    23 => '0' & "000000" &  '0' & x"00800000",
    24 => '0' & "000000" &  '0' & x"01000000",
    25 => '0' & "000000" &  '0' & x"02000000",
    26 => '0' & "000000" &  '0' & x"04000000",
    27 => '0' & "000000" &  '0' & x"08000000",
    28 => '0' & "000000" &  '0' & x"10000000",
    29 => '0' & "000000" &  '0' & x"20000000",
    30 => '0' & "000000" &  '0' & x"40000000",
    31 => '0' & "000000" &  '0' & x"80000000",
    32 => '0' & "000000" &  '1' & x"00000000",
    33 => '1' & "000000" &  '0' & x"00000000",
    34 => '0' & "000000" &  '0' & x"00000000",
    35 => '0' & "000000" &  '0' & x"00000000",
    36 => '0' & "000000" &  '0' & x"00000000",
    37 => '0' & "000000" &  '0' & x"00000000",
    38 => '0' & "000000" &  '0' & x"00000000",
    39 => '0' & "000000" &  '0' & x"00000000",
    40 => '0' & "000000" &  '0' & x"00000000",
    41 => '0' & "000000" &  '0' & x"00000000",
    42 => '0' & "000000" &  '0' & x"00000000",
    43 => '0' & "000000" &  '0' & x"00000000",
    44 => '0' & "000000" &  '0' & x"00000000",
    45 => '0' & "000000" &  '0' & x"00000000",
    46 => '0' & "000000" &  '0' & x"00000000",
    47 => '0' & "000000" &  '0' & x"00000000",
    48 => '0' & "000000" &  '0' & x"00000000",
    49 => '0' & "000000" &  '0' & x"00000000",
    50 => '0' & "000000" &  '0' & x"00000000",
    51 => '0' & "000000" &  '0' & x"00000000",
    52 => '0' & "000000" &  '0' & x"00000000",
    53 => '0' & "000000" &  '0' & x"00000000",
    54 => '0' & "000000" &  '0' & x"00000000",
    55 => '0' & "000000" &  '0' & x"00000000",
    56 => '0' & "000000" &  '0' & x"00000000",
    57 => '0' & "000000" &  '0' & x"00000000",
    58 => '0' & "000000" &  '0' & x"00000000",
    59 => '0' & "000000" &  '0' & x"00000000",
    60 => '0' & "000000" &  '0' & x"00000000",
    61 => '0' & "000000" &  '0' & x"00000000",
    62 => '0' & "000000" &  '0' & x"00000000",
    63 => '0' & "000000" &  '0' & x"00000000",
    64 => '0' & "000000" &  '0' & x"00000000",
    65 => '0' & "000000" &  '0' & x"00000000",
    66 => '0' & "000000" &  '0' & x"00000000",
    67 => '0' & "000000" &  '0' & x"00000000",
    68 => '0' & "000000" &  '0' & x"00000000",
    69 => '0' & "000000" &  '0' & x"00000000",
    70 => '0' & "000000" &  '0' & x"00000000",
    71 => '0' & "000000" &  '0' & x"00000000",
    72 => '0' & "000000" &  '0' & x"00000000",
    73 => '0' & "000000" &  '0' & x"00000000",
    74 => '0' & "000000" &  '0' & x"00000000",
    75 => '0' & "000000" &  '0' & x"00000000",
    76 => '0' & "000000" &  '0' & x"00000000",
    77 => '0' & "000000" &  '0' & x"00000000",
    78 => '0' & "000000" &  '0' & x"00000000",
    79 => '0' & "000000" &  '0' & x"00000000",
    80 => '0' & "000000" &  '0' & x"00000000",
    81 => '0' & "000000" &  '0' & x"00000000",
    82 => '0' & "000000" &  '0' & x"00000000",
    83 => '0' & "000000" &  '0' & x"00000000",
    84 => '0' & "000000" &  '0' & x"00000000",
    85 => '0' & "000000" &  '0' & x"00000000",
    86 => '0' & "000000" &  '0' & x"00000000",
    87 => '0' & "000000" &  '0' & x"00000000",
    88 => '0' & "000000" &  '0' & x"00000000",
    89 => '0' & "000000" &  '0' & x"00000000",
    90 => '0' & "000000" &  '0' & x"00000000",
    91 => '0' & "000000" &  '0' & x"00000000",
    92 => '0' & "000000" &  '0' & x"00000000",
    93 => '0' & "000000" &  '0' & x"00000000",
    94 => '0' & "000000" &  '0' & x"00000000",
    95 => '0' & "000000" &  '0' & x"00000000",
    96 => '0' & "000000" &  '0' & x"00000000",
    97 => '0' & "000000" &  '0' & x"00000000",
    98 => '0' & "000000" &  '0' & x"00000000",
    99 => '0' & "000000" &  '0' & x"00000000",
    100 => '0' & "000000" &  '0' & x"00000000",
    101 => '0' & "000000" &  '0' & x"00000000",
    102 => '0' & "000000" &  '0' & x"00000000",
    103 => '0' & "000000" &  '0' & x"00000000",
    104 => '0' & "000000" &  '0' & x"00000000",
    105 => '0' & "000000" &  '0' & x"00000000",
    106 => '0' & "000000" &  '0' & x"00000000",
    107 => '0' & "000000" &  '0' & x"00000000",
    108 => '0' & "000000" &  '0' & x"00000000",
    109 => '0' & "000000" &  '0' & x"00000000",
    110 => '0' & "000000" &  '0' & x"00000000",
    111 => '0' & "000000" &  '0' & x"00000000",
    112 => '0' & "000000" &  '0' & x"00000000",
    113 => '0' & "000000" &  '0' & x"00000000",
    114 => '0' & "000000" &  '0' & x"00000000",
    115 => '0' & "000000" &  '0' & x"00000000",
    116 => '0' & "000000" &  '0' & x"00000000",
    117 => '0' & "000000" &  '0' & x"00000000",
    118 => '0' & "000000" &  '0' & x"00000000",
    119 => '0' & "000000" &  '0' & x"00000000",
    120 => '0' & "000000" &  '0' & x"00000000",
    121 => '1' & "000000" &  '0' & x"00000000",
    122 => '1' & "000000" &  '0' & x"00000000",
    123 => '1' & "000000" &  '0' & x"00000000",
    124 => '1' & "000000" &  '0' & x"00000000",
    125 => '0' & "000001" &  '0' & x"00000000",
    126 => '0' & "000010" &  '0' & x"00000000",
    127 => '0' & "000011" &  '0' & x"00000000",
    128 => '0' & "000100" &  '0' & x"00000000",
    129 => '0' & "000101" &  '0' & x"00000000",
    130 => '0' & "000110" &  '0' & x"00000000",
    131 => '0' & "000111" &  '0' & x"00000000",
    132 => '0' & "001000" &  '0' & x"00000000",
    133 => '0' & "001001" &  '0' & x"00000000",
    134 => '0' & "001010" &  '0' & x"00000000",
    135 => '0' & "001011" &  '0' & x"00000000",
    136 => '0' & "001100" &  '0' & x"00000000",
    137 => '0' & "001101" &  '0' & x"00000000",
    138 => '0' & "001110" &  '0' & x"00000000",
    139 => '0' & "001111" &  '0' & x"00000000",
    140 => '0' & "010000" &  '0' & x"00000000",
    141 => '0' & "010001" &  '0' & x"00000000",
    142 => '0' & "010010" &  '0' & x"00000000",
    143 => '0' & "010011" &  '0' & x"00000000",
    144 => '0' & "010100" &  '0' & x"00000000",
    145 => '0' & "010101" &  '0' & x"00000000",
    146 => '0' & "010110" &  '0' & x"00000000",
    147 => '0' & "010111" &  '0' & x"00000000",
    148 => '0' & "011000" &  '0' & x"00000000",
    149 => '0' & "011001" &  '0' & x"00000000",
    150 => '0' & "011010" &  '0' & x"00000000",
    151 => '0' & "011011" &  '0' & x"00000000",
    152 => '0' & "011100" &  '0' & x"00000000",
    153 => '0' & "011101" &  '0' & x"00000000",
    154 => '0' & "011110" &  '0' & x"00000000",
    155 => '0' & "011111" &  '0' & x"00000000",
    156 => '0' & "100000" &  '0' & x"00000000",
    157 => '0' & "100001" &  '0' & x"00000000",
    158 => '0' & "100010" &  '0' & x"00000000",
    159 => '0' & "000000" &  '0' & x"00000000",
    160 => '0' & "000000" &  '0' & x"00000000",
    161 => '0' & "000000" &  '0' & x"00000000",
    162 => '0' & "000000" &  '0' & x"00000000",
    163 => '0' & "000000" &  '0' & x"00000000",
    164 => '0' & "000000" &  '0' & x"00000000",
    165 => '0' & "000000" &  '0' & x"00000000",
    166 => '0' & "000000" &  '0' & x"00000000",
    167 => '0' & "000000" &  '0' & x"00000000",
    168 => '0' & "000000" &  '0' & x"00000000",
    169 => '0' & "000000" &  '0' & x"00000000",
    170 => '0' & "000000" &  '0' & x"00000000",
    171 => '0' & "000000" &  '0' & x"00000000",
    172 => '0' & "000000" &  '0' & x"00000000",
    173 => '0' & "000000" &  '0' & x"00000000",
    174 => '0' & "000000" &  '0' & x"00000000",
    175 => '0' & "000000" &  '0' & x"00000000",
    176 => '0' & "000000" &  '0' & x"00000000",
    177 => '0' & "000000" &  '0' & x"00000000",
    178 => '0' & "000000" &  '0' & x"00000000",
    179 => '0' & "000000" &  '0' & x"00000000",
    180 => '0' & "000000" &  '0' & x"00000000",
    181 => '0' & "000000" &  '0' & x"00000000",
    182 => '0' & "000000" &  '0' & x"00000000",
    183 => '0' & "000000" &  '0' & x"00000000",
    184 => '0' & "000000" &  '0' & x"00000000",
    185 => '0' & "000000" &  '0' & x"00000000",
    186 => '0' & "000000" &  '0' & x"00000000",
    187 => '0' & "000000" &  '0' & x"00000000",
    188 => '0' & "000000" &  '0' & x"00000000",
    189 => '0' & "000000" &  '0' & x"00000000",
    190 => '0' & "000000" &  '0' & x"00000000",
    191 => '0' & "000000" &  '0' & x"00000000",
    192 => '0' & "000000" &  '0' & x"00000000",
    193 => '0' & "000000" &  '0' & x"00000000",
    194 => '0' & "000000" &  '0' & x"00000000",
    195 => '0' & "000000" &  '0' & x"00000000",
    196 => '0' & "000000" &  '0' & x"00000000",
    197 => '0' & "000000" &  '0' & x"00000000",
    198 => '0' & "000000" &  '0' & x"00000000",
    199 => '0' & "000000" &  '0' & x"00000000",
    200 => '0' & "000000" &  '0' & x"00000000",
    201 => '0' & "000000" &  '0' & x"00000000",
    202 => '0' & "000000" &  '0' & x"00000000",
    203 => '0' & "000000" &  '0' & x"00000000",
    204 => '0' & "000000" &  '0' & x"00000000",
    205 => '0' & "000000" &  '0' & x"00000000",
    206 => '0' & "000000" &  '0' & x"00000000",
    207 => '0' & "000000" &  '0' & x"00000000",
    208 => '0' & "000000" &  '0' & x"00000000",
    209 => '0' & "000000" &  '0' & x"00000000",
    210 => '0' & "000000" &  '0' & x"00000000",
    211 => '0' & "000000" &  '0' & x"00000000",
    212 => '0' & "000000" &  '0' & x"00000000",
    213 => '0' & "000000" &  '0' & x"00000000",
    214 => '0' & "000000" &  '0' & x"00000000",
    215 => '0' & "000000" &  '0' & x"00000000",
    216 => '0' & "000000" &  '0' & x"00000000",
    217 => '0' & "000000" &  '0' & x"00000000",
    218 => '0' & "000000" &  '0' & x"00000000",
    219 => '0' & "000000" &  '0' & x"00000000",
    220 => '0' & "000000" &  '0' & x"00000000",
    221 => '0' & "000000" &  '0' & x"00000000",
    222 => '0' & "000000" &  '0' & x"00000000",
    223 => '0' & "000000" &  '0' & x"00000000",
    224 => '0' & "000000" &  '0' & x"00000000",
    225 => '0' & "000000" &  '0' & x"00000000",
    226 => '0' & "000000" &  '0' & x"00000000",
    227 => '0' & "000000" &  '0' & x"00000000",
    228 => '0' & "000000" &  '0' & x"00000000",
    229 => '0' & "000000" &  '0' & x"00000000",
    230 => '0' & "000000" &  '0' & x"00000000",
    231 => '0' & "000000" &  '0' & x"00000000",
    232 => '0' & "000000" &  '0' & x"00000000",
    233 => '0' & "000000" &  '0' & x"00000000",
    234 => '0' & "000000" &  '0' & x"00000000",
    235 => '0' & "000000" &  '0' & x"00000000",
    236 => '0' & "000000" &  '0' & x"00000000",
    237 => '0' & "000000" &  '0' & x"00000000",
    238 => '0' & "000000" &  '0' & x"00000000",
    239 => '0' & "000000" &  '0' & x"00000000",
    240 => '0' & "000000" &  '0' & x"00000000",
    241 => '0' & "000000" &  '0' & x"00000000",
    242 => '0' & "000000" &  '0' & x"00000000",
    243 => '0' & "000000" &  '0' & x"00000000",
    244 => '0' & "000000" &  '0' & x"00000000",
    245 => '0' & "000000" &  '0' & x"00000000",
    246 => '0' & "000000" &  '0' & x"00000000",
    247 => '0' & "000000" &  '0' & x"00000000",
    248 => '0' & "000000" &  '0' & x"00000000",
    249 => '0' & "000000" &  '0' & x"00000000",
    250 => '1' & "000000" &  '0' & x"00000000",
    251 => '1' & "000000" &  '0' & x"00000000",
    252 => '1' & "000000" &  '0' & x"00000000",
    253 => '1' & "000000" &  '0' & x"00000000",
    254 => '0' & "000000" &  '0' & x"00000000",
    255 => '1' & "000000" &  '0' & x"00000000"
    );

end package;
