----------------------------------------------------------------------------------
-- Company: DHBW
-- Engineer: Levi Bohnacker
-- 
-- Create Date: 05/23/2021 11:12:41 AM
-- Design Name: CSR_top
-- Module Name: sim_CSR_top_UV_2_pkg
-- Project Name: EDRICO
-- Target Devices: Arty Z7
-- Tool Versions: 
-- Description: 
--  this package contains stimuli and verification dat for the 
--  sim_CSR_top_UV_2_tb.vhd testbench.
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


----------------------------------------------------------------------------------
--PACKAGE
----------------------------------------------------------------------------------
package sim_CSR_top_UV_2_pkg is 
----------------------------------------------------------------------------------
--types
----------------------------------------------------------------------------------
---stimulation dat
--control_stim(13) = CSR_write, control_stim(12) = CSR_read, control_stim(11 downto 0) = CSR_address
type control_stim is array(natural range <>) of std_logic_vector(13 downto 0);
type data_stim is array(natural range  <>) of std_logic_vector(31 downto 0);
--input_stim(2) = MSIP_dra, input_stim(1) = MTIP_dra, input_stim(0) = instr_finished
type input_stim  is array(natural range <>) of std_logic_vector(2 downto 0);

--verification data
--result_vect(32) = illegal_instruction_exception, result_vect(31 downto 0) = data_out
type result_vect is array(natural range <>) of std_logic_vector(32 downto 0);

----------------------------------------------------------------------------------
--constants
----------------------------------------------------------------------------------
constant results : result_vect(255 downto 0) :=
    (
    0 => '0' & x"00000000", 
    1 => '0' & x"00000000", 
    2 => '0' & x"00000000", 
    3 => '0' & x"00000000", 
    4 => '0' & x"00000000", 
    5 => '0' & x"00000000", 
    6 => '0' & x"00000000", 
    7 => '0' & x"00000000", 
    8 => '0' & x"00000000", 
    9 => '0' & x"00000000", 
    10 => '0' & x"00000000", 
    11 => '0' & x"00000000", 
    12 => '0' & x"00000000", 
    13 => '0' & x"00000000", 
    14 => '0' & x"00000000", 
    15 => '0' & x"00000000", 
    16 => '0' & x"00000000", 
    17 => '0' & x"00000000", 
    18 => '0' & x"00000000", 
    19 => '0' & x"00000000", 
    20 => '0' & x"00000000", 
    21 => '0' & x"00000000", 
    22 => '0' & x"00000000", 
    23 => '0' & x"00000000", 
    24 => '0' & x"00000000", 
    25 => '0' & x"00000000", 
    26 => '0' & x"00000000", 
    27 => '0' & x"00000000", 
    28 => '0' & x"00000000", 
    29 => '0' & x"00000000", 
    30 => '0' & x"00000000", 
    31 => '0' & x"00000000", 
    32 => '0' & x"00000000", 
    33 => '0' & x"00000000", 
    34 => '1' & x"00000000", 
    35 => '0' & x"00000000", 
    36 => '0' & x"00000000", 
    37 => '0' & x"00000000", 
    38 => '0' & x"00000000", 
    39 => '0' & x"00000000", 
    40 => '0' & x"00000000", 
    41 => '0' & x"00000000", 
    42 => '0' & x"00000000", 
    43 => '0' & x"00000000", 
    44 => '0' & x"00000000", 
    45 => '0' & x"00000000", 
    46 => '0' & x"00000000", 
    47 => '0' & x"00000000", 
    48 => '0' & x"00000000", 
    49 => '0' & x"00000000", 
    50 => '0' & x"00000000", 
    51 => '0' & x"00000000", 
    52 => '0' & x"00000000", 
    53 => '0' & x"00000000", 
    54 => '0' & x"00000000", 
    55 => '0' & x"00000000", 
    56 => '0' & x"00000000", 
    57 => '0' & x"00000000", 
    58 => '0' & x"00000000", 
    59 => '0' & x"00000000", 
    60 => '0' & x"00000000", 
    61 => '0' & x"00000000", 
    62 => '0' & x"00000000", 
    63 => '0' & x"00000000", 
    64 => '0' & x"00000000", 
    65 => '0' & x"00000000", 
    66 => '0' & x"00000000", 
    67 => '0' & x"00000000", 
    68 => '0' & x"00000000", 
    69 => '0' & x"00000000", 
    70 => '0' & x"00000000", 
    71 => '0' & x"00000000", 
    72 => '0' & x"00000000", 
    73 => '0' & x"00000000", 
    74 => '0' & x"00000000", 
    75 => '0' & x"00000000", 
    76 => '0' & x"00000000", 
    77 => '0' & x"00000000", 
    78 => '0' & x"00000000", 
    79 => '0' & x"00000000", 
    80 => '0' & x"00000000", 
    81 => '0' & x"00000000", 
    82 => '0' & x"00000000", 
    83 => '0' & x"00000000", 
    84 => '0' & x"00000000", 
    85 => '0' & x"00000000", 
    86 => '0' & x"00000000", 
    87 => '0' & x"00000000", 
    88 => '0' & x"00000000", 
    89 => '0' & x"00000000", 
    90 => '0' & x"00000000", 
    91 => '0' & x"00000000", 
    92 => '0' & x"00000000", 
    93 => '0' & x"00000000", 
    94 => '0' & x"00000000", 
    95 => '0' & x"00000000", 
    96 => '0' & x"00000000", 
    97 => '0' & x"00000000", 
    98 => '0' & x"00000000", 
    99 => '0' & x"00000000", 
    100 => '0' & x"00000000", 
    101 => '0' & x"00000000", 
    102 => '0' & x"00000000", 
    103 => '0' & x"00000000", 
    104 => '0' & x"00000000", 
    105 => '0' & x"00000000", 
    106 => '0' & x"00000000", 
    107 => '0' & x"00000000", 
    108 => '0' & x"00000000", 
    109 => '0' & x"00000000", 
    110 => '0' & x"00000000", 
    111 => '0' & x"00000000", 
    112 => '0' & x"00000000", 
    113 => '0' & x"00000000", 
    114 => '0' & x"00000000", 
    115 => '0' & x"00000000", 
    116 => '0' & x"00000000", 
    117 => '0' & x"00000000", 
    118 => '0' & x"00000000", 
    119 => '0' & x"00000000", 
    120 => '0' & x"00000000", 
    121 => '0' & x"00000000", 
    122 => '1' & x"00000000", 
    123 => '1' & x"00000000", 
    124 => '1' & x"00000000", 
    125 => '1' & x"00000000", 
    126 => '0' & x"00001808", --mstatus
    127 => '0' & x"FFFFFFFF", --minstretH
    128 => '0' & x"00000088", --mie
    129 => '0' & x"0A000000", --mtvec
    130 => '0' & x"00000000", --mcountinhibit
    131 => '0' & x"DEADAFFE", --mscratch
    132 => '0' & x"00037512", --mepc
    133 => '0' & x"BADC0DED", --mcause
    134 => '0' & x"ABBABABA", --mtval
    135 => '0' & x"00000088", --mip
    136 => '0' & "10000000" & "10011001" & "10011111" & "10001101", --pmpcfg0
    137 => '0' & "10011011" & "10011011" & "10011011" & "10001011", --pmpcfg1
    138 => '0' & "10001111" & "10000000" & "10010011" & "10011000", --pmpcfg2
    139 => '0' & "10000101" & "10000101" & "10000101" & "10011111", --pmpcfg3
    140 => '0' & x"00400000", --pmpaddr0
    141 => '0' & x"005FFFFF", --pmpaddr1
    142 => '0' & x"009FFFFF", --pmpaddr2
    143 => '0' & x"00C00000", --pmpaddr3
    144 => '0' & x"14000000", --pmpaddr4
    145 => '0' & x"1400001F", --pmpaddr5
    146 => '0' & x"1400005F", --pmpaddr6
    147 => '0' & x"1400009F", --pmpaddr7
    148 => '0' & x"140000DF", --pmpaddr8
    149 => '0' & x"14000100", --pmpaddr9
    150 => '0' & x"14000100", --pmpaddr10
    151 => '0' & x"FFFFFFFF", --pmpaddr11
    152 => '0' & x"009FFFFF", --pmpaddr12
    153 => '0' & x"005FFFFF", --pmpaddr13
    154 => '0' & x"003FFFFF", --pmpaddr14
    155 => '0' & x"003FFFFF", --pmpaddr15
    156 => '0' & x"10000096", --mcycle
    157 => '0' & x"10000013", --minstret
    158 => '0' & x"FFFFFFFF", --mcycleH
    159 => '0' & x"00000100", --misa
    160 => '0' & x"00000000", 
    161 => '0' & x"00000000", 
    162 => '0' & x"00000000", 
    163 => '0' & x"00000000", 
    164 => '0' & x"00000000", 
    165 => '0' & x"00000000", 
    166 => '0' & x"00000000", 
    167 => '0' & x"00000000", 
    168 => '0' & x"00000000", 
    169 => '0' & x"00000000", 
    170 => '0' & x"00000000", 
    171 => '0' & x"00000000", 
    172 => '0' & x"00000000", 
    173 => '0' & x"00000000", 
    174 => '0' & x"00000000", 
    175 => '0' & x"00000000", 
    176 => '0' & x"00000000", 
    177 => '0' & x"00000000", 
    178 => '0' & x"00000000", 
    179 => '0' & x"00000000", 
    180 => '0' & x"00000000", 
    181 => '0' & x"00000000", 
    182 => '0' & x"00000000", 
    183 => '0' & x"00000000", 
    184 => '0' & x"00000000", 
    185 => '0' & x"00000000", 
    186 => '0' & x"00000000", 
    187 => '0' & x"00000000", 
    188 => '0' & x"00000000", 
    189 => '0' & x"00000000", 
    190 => '0' & x"00000000", 
    191 => '0' & x"00000000", 
    192 => '0' & x"00000000", 
    193 => '0' & x"00000000", 
    194 => '0' & x"00000000", 
    195 => '0' & x"00000000", 
    196 => '0' & x"00000000", 
    197 => '0' & x"00000000", 
    198 => '0' & x"00000000", 
    199 => '0' & x"00000000", 
    200 => '0' & x"00000000", 
    201 => '0' & x"00000000", 
    202 => '0' & x"00000000", 
    203 => '0' & x"00000000", 
    204 => '0' & x"00000000", 
    205 => '0' & x"00000000", 
    206 => '0' & x"00000000", 
    207 => '0' & x"00000000", 
    208 => '0' & x"00000000", 
    209 => '0' & x"00000000", 
    210 => '0' & x"00000000", 
    211 => '0' & x"00000000", 
    212 => '0' & x"00000000", 
    213 => '0' & x"00000000", 
    214 => '0' & x"00000000", 
    215 => '0' & x"00000000", 
    216 => '0' & x"00000000", 
    217 => '0' & x"00000000", 
    218 => '0' & x"00000000", 
    219 => '0' & x"00000000", 
    220 => '0' & x"00000000", 
    221 => '0' & x"00000000", 
    222 => '0' & x"00000000", 
    223 => '0' & x"00000000", 
    224 => '0' & x"00000000", 
    225 => '0' & x"00000000", 
    226 => '0' & x"00000000", 
    227 => '0' & x"00000000", 
    228 => '0' & x"00000000", 
    229 => '0' & x"00000000", 
    230 => '0' & x"00000000", 
    231 => '0' & x"00000000", 
    232 => '0' & x"00000000", 
    233 => '0' & x"00000000", 
    234 => '0' & x"00000000", 
    235 => '0' & x"00000000", 
    236 => '0' & x"00000000", 
    237 => '0' & x"00000000", 
    238 => '0' & x"00000000", 
    239 => '0' & x"00000000", 
    240 => '0' & x"00000000", 
    241 => '0' & x"00000000", 
    242 => '0' & x"00000000", 
    243 => '0' & x"00000000", 
    244 => '0' & x"00000000", 
    245 => '0' & x"00000000", 
    246 => '0' & x"00000000", 
    247 => '0' & x"00000000", 
    248 => '0' & x"00000000", 
    249 => '0' & x"00000000", 
    250 => '0' & x"00000000", 
    251 => '1' & x"00000000", --faulty address
    252 => '1' & x"00000000", --faulty address
    253 => '1' & x"00000000", --faulty address
    254 => '1' & x"00000000", --faulty address
    255 => '0' & x"00000000" --faulty address
    );

--input_stim(2) = MSIP_dra, input_stim(1) = MTIP_dra, input_stim(0) = instr_finished
constant stimulus_input : input_stim(7 downto 0) :=
    (
    0 => "000",
    1 => "000",
    2 => "000",
    3 => "000",
    4 => "110",
    5 => "110",
    6 => "110",
    7 => "111"
    );

constant stimulus_data : data_stim(255 downto 0) :=
    (
    0 => x"00000005",   --disable cy and ir counter
    1 => x"10000000",   --starting value for mcycle:    0xFFFFFFFF10000000
    2 => x"FFFFFFFF", 
    3 => x"10000000",   --starting value for minstret:  0xFFFFFFFF10000000
    4 => x"FFFFFFFF",
    5 => x"00000000",   --activate cy and ir counter
    6 => x"00000008",   --set MIE and clear MPIE in mstatus
    7 => x"00000088",   --enable mtip and msip interrupts => should be high
    8 => x"00000000",   --clear mtip and msip bit
    9 => x"0A000000",   --mtvec (base address = 0x0A000000, mode: direct)
    10 => x"DEADAFFE",  --dummy data to mscratch
    11 => x"00037512",  --dummy data to mepc
    12 => x"BADC0DED",  --dummy data to mcause
    13 => x"ABBABABA",   --dummy data to mtval
    --pmpregister config same as in sim_PMP_checker_UV_2
    14 => "10000000" & "10011001" & "10011111" & "10001101",
    15 => "10011011" & "10011011" & "10011011" & "10001011",
    16 => "10001111" & "10000000" & "10010011" & "10011000",
    17 => "10000101" & "10000101" & "10000101" & "10011111",
    18 => x"00400000",  --ROM0
    19 => x"005FFFFF",  --RAM0
    20 => x"009FFFFF",  --ROM1
    21 => x"00C00000",  --RAM1_L
    22 => x"14000000",  --RAM1
    23 => x"1400001F",  --RAM2
    24 => x"1400005F",  --RAM3
    25 => x"1400009F",  --RAM4
    26 => x"140000DF",  --Region0
    27 => x"14000100",  --Region1
    28 => x"14000100",  --Region2_L
    29 => x"FFFFFFFF",  --Region2
    30 => x"009FFFFF",  --ROM1 redefind
    31 => x"005FFFFF",  --not used
    32 => x"003FFFFF",  --not used
    33 => x"003FFFFF",  --not used
    34 => x"10293812",  --dummy data to misa
    --random generated data for read, read-only registers and error tests
    35	=> x"F768DD4F",	--mhpmevent3
    36	=> x"D3695828",	--mhpmevent4
    37	=> x"C824EC0F",	--mhpmevent5
    38	=> x"83A96D7A",	--mhpmevent6
    39	=> x"064649F8",	--mhpmevent7
    40	=> x"C9E29349",	--mhpmevent8
    41	=> x"D4839B5F",	--mhpmevent9
    42	=> x"4DF8952B",	--mhpmevent10
    43	=> x"45787E34",	--mhpmevent11
    44	=> x"B39CD499",	--mhpmevent12
    45	=> x"C26B4139",	--mhpmevent13
    46	=> x"0A821692",	--mhpmevent14
    47	=> x"65301D89",	--mhpmevent15
    48	=> x"3F5FAF76",	--mhpmevent16
    49	=> x"60EA493A",	--mhpmevent17
    50	=> x"855B52DA",	--mhpmevent18
    51	=> x"0FFEC211",	--mhpmevent19
    52	=> x"00D2BC79",	--mhpmevent20
    53	=> x"5A2FCA27",	--mhpmevent21
    54	=> x"EAC7BDF3",	--mhpmevent22
    55	=> x"9778F9EF",	--mhpmevent23
    56	=> x"E0DA471B",	--mhpmevent24
    57	=> x"468DEEE1",	--mhpmevent25
    58	=> x"6250095D",	--mhpmevent26
    59	=> x"680F3C7F",	--mhpmevent27
    60	=> x"2B2A452B",	--mhpmevent28
    61	=> x"5220A144",	--mhpmevent29
    62	=> x"187773FB",	--mhpmevent30
    63	=> x"F31D575D",	--mhpmevent31
    64	=> x"B7F9232C",	--mhpmcounter3
    65	=> x"08CB99D6",	--mhpmcounter4
    66	=> x"6B6BDB15",	--mhpmcounter5
    67	=> x"346AF93D",	--mhpmcounter6
    68	=> x"7ECF6E71",	--mhpmcounter7
    69	=> x"6F4224BB",	--mhpmcounter8
    70	=> x"F2C52B27",	--mhpmcounter9
    71	=> x"3892790C",	--mhpmcounter10
    72	=> x"992BFC92",	--mhpmcounter11
    73	=> x"3CA3F55D",	--mhpmcounter12
    74	=> x"C0FB35F7",	--mhpmcounter13
    75	=> x"4C29AA71",	--mhpmcounter14
    76	=> x"51EF5C53",	--mhpmcounter15
    77	=> x"77D586B8",	--mhpmcounter16
    78	=> x"62CEAFEC",	--mhpmcounter17
    79	=> x"FC838594",	--mhpmcounter18
    80	=> x"458B978E",	--mhpmcounter19
    81	=> x"67EA468E",	--mhpmcounter20
    82	=> x"0DD51DE1",	--mhpmcounter21
    83	=> x"B54F6C16",	--mhpmcounter22
    84	=> x"34017B84",	--mhpmcounter23
    85	=> x"8FA88CD5",	--mhpmcounter24
    86	=> x"EDAAD6FE",	--mhpmcounter25
    87	=> x"6F1BDBE2",	--mhpmcounter26
    88	=> x"E59A5B7F",	--mhpmcounter27
    89	=> x"DE53ECD4",	--mhpmcounter28
    90	=> x"A44613A4",	--mhpmcounter29
    91	=> x"2847D97C",	--mhpmcounter30
    92	=> x"DEFDDA4B",	--mhpmcounter31
    93	=> x"5977391C",	--mhpmcounterH3
    94	=> x"CDF9CB42",	--mhpmcounterH4
    95	=> x"E40CFC9D",	--mhpmcounterH5
    96	=> x"07C1058D",	--mhpmcounterH6
    97	=> x"11742DAC",	--mhpmcounterH7
    98	=> x"005CBE88",	--mhpmcounterH8
    99	=> x"82DCC624",	--mhpmcounterH9
    100	=> x"7F3DBED8",	--mhpmcounterH10
    101	=> x"F3AA61E0",	--mhpmcounterH11
    102	=> x"83B5168D",	--mhpmcounterH12
    103	=> x"B213DDCE",	--mhpmcounterH13
    104	=> x"901D115A",	--mhpmcounterH14
    105	=> x"6C5E650E",	--mhpmcounterH15
    106	=> x"91AD4AD2",	--mhpmcounterH16
    107	=> x"C4B5A292",	--mhpmcounterH17
    108	=> x"EADD9A59",	--mhpmcounterH18
    109	=> x"78CF9580",	--mhpmcounterH19
    110	=> x"858CBCDF",	--mhpmcounterH20
    111	=> x"D4A102B8",	--mhpmcounterH21
    112	=> x"4BF4E08B",	--mhpmcounterH22
    113	=> x"F5319334",	--mhpmcounterH23
    114	=> x"E9FB5B9C",	--mhpmcounterH24
    115	=> x"72E45486",	--mhpmcounterH25
    116	=> x"D6E86335",	--mhpmcounterH26
    117	=> x"8A904213",	--mhpmcounterH27
    118	=> x"ABD39E66",	--mhpmcounterH28
    119	=> x"2581B17A",	--mhpmcounterH29
    120	=> x"C2A5CEA0",	--mhpmcounterH30
    121	=> x"ED171E93",	--mhpmcounterH31
    122	=> x"1FFCB24E",	--mvendorid
    123	=> x"5DE0DAE1",	--marchid
    124	=> x"CB45BE1E",	--mimpid
    125	=> x"4438FDBA",	--mhartid
    126	=> x"4FEF482A",	--mstatus
    127	=> x"BE8D2C89",	--minstretH
    128	=> x"741A2A88",	--mie
    129	=> x"7736F91A",	--mtvec
    130	=> x"B7E1A78C",	--mcountinhibit
    131	=> x"57DD978E",	--mscratch
    132	=> x"5369A92A",	--mepc
    133	=> x"B63E86A8",	--mcause
    134	=> x"3B5B5C69",	--mtval
    135	=> x"C8266287",	--mip
    136	=> x"3E65D9F8",	--pmpcfg0
    137	=> x"3026FAB1",	--pmpcfg1
    138	=> x"091DFF87",	--pmpcfg2
    139	=> x"BE5FD367",	--pmpcfg3
    140	=> x"57816037",	--pmpaddr0
    141	=> x"76D616AA",	--pmpaddr1
    142	=> x"389FC79E",	--pmpaddr2
    143	=> x"273AEDB5",	--pmpaddr3
    144	=> x"F9BA11B3",	--pmpaddr4
    145	=> x"471E06AB",	--pmpaddr5
    146	=> x"36B95DFD",	--pmpaddr6
    147	=> x"2D6275E8",	--pmpaddr7
    148	=> x"0BF81BF4",	--pmpaddr8
    149	=> x"9C3B87DA",	--pmpaddr9
    150	=> x"EC02A8B3",	--pmpaddr10
    151	=> x"1A8B5101",	--pmpaddr11
    152	=> x"4F96BBBE",	--pmpaddr12
    153	=> x"3DB32D9C",	--pmpaddr13
    154	=> x"606C339F",	--pmpaddr14
    155	=> x"089449EE",	--pmpaddr15
    156	=> x"422B16C9",	--mcycle
    157	=> x"D3733D28",	--minstret
    158	=> x"E809945D",	--mcycleH
    159	=> x"9A84FA24",	--misa
    160	=> x"42E56EFA",	--mhpmevent3
    161	=> x"75A38D61",	--mhpmevent4
    162	=> x"E0031CAD",	--mhpmevent5
    163	=> x"9B1425C4",	--mhpmevent6
    164	=> x"87A11777",	--mhpmevent7
    165	=> x"E6A99911",	--mhpmevent8
    166	=> x"4727E3DD",	--mhpmevent9
    167	=> x"97F1A9CE",	--mhpmevent10
    168	=> x"DF78A236",	--mhpmevent11
    169	=> x"62590BE8",	--mhpmevent12
    170	=> x"6B24E006",	--mhpmevent13
    171	=> x"0A203301",	--mhpmevent14
    172	=> x"3FE249D6",	--mhpmevent15
    173	=> x"5D6F1353",	--mhpmevent16
    174	=> x"5D82AD7C",	--mhpmevent17
    175	=> x"199715CE",	--mhpmevent18
    176	=> x"EA8C288A",	--mhpmevent19
    177	=> x"8476D963",	--mhpmevent20
    178	=> x"ECD7BB54",	--mhpmevent21
    179	=> x"9FD713C8",	--mhpmevent22
    180	=> x"A78E9B58",	--mhpmevent23
    181	=> x"E09A2F97",	--mhpmevent24
    182	=> x"1693EA9D",	--mhpmevent25
    183	=> x"4BA40930",	--mhpmevent26
    184	=> x"5F8FC0EB",	--mhpmevent27
    185	=> x"77E62B61",	--mhpmevent28
    186	=> x"443E550E",	--mhpmevent29
    187	=> x"F7B1D476",	--mhpmevent30
    188	=> x"7021AECE",	--mhpmevent31
    189	=> x"D2C2C0E4",	--mhpmcounter3
    190	=> x"0290D1C7",	--mhpmcounter4
    191	=> x"ACBF21AE",	--mhpmcounter5
    192	=> x"6FEBE101",	--mhpmcounter6
    193	=> x"4416FE63",	--mhpmcounter7
    194	=> x"1C3607D3",	--mhpmcounter8
    195	=> x"12354CB0",	--mhpmcounter9
    196	=> x"823D35F0",	--mhpmcounter10
    197	=> x"AD5F67B7",	--mhpmcounter11
    198	=> x"C58DD517",	--mhpmcounter12
    199	=> x"4E669940",	--mhpmcounter13
    200	=> x"CE564CFF",	--mhpmcounter14
    201	=> x"AADB5344",	--mhpmcounter15
    202	=> x"CB43106C",	--mhpmcounter16
    203	=> x"82C01AB2",	--mhpmcounter17
    204	=> x"467D1136",	--mhpmcounter18
    205	=> x"99790019",	--mhpmcounter19
    206	=> x"C68CB3FE",	--mhpmcounter20
    207	=> x"D0B9FE13",	--mhpmcounter21
    208	=> x"93FE87A9",	--mhpmcounter22
    209	=> x"F5EABC1F",	--mhpmcounter23
    210	=> x"E0B6B205",	--mhpmcounter24
    211	=> x"C83BF2FF",	--mhpmcounter25
    212	=> x"A88E534A",	--mhpmcounter26
    213	=> x"A2569FB9",	--mhpmcounter27
    214	=> x"CEB7E3CD",	--mhpmcounter28
    215	=> x"E40149D3",	--mhpmcounter29
    216	=> x"B48C01BB",	--mhpmcounter30
    217	=> x"52EBADD4",	--mhpmcounter31
    218	=> x"74BE5E63",	--mhpmcounterH3
    219	=> x"0332BF1B",	--mhpmcounterH4
    220	=> x"91C387D3",	--mhpmcounterH5
    221	=> x"C9B9F38C",	--mhpmcounterH6
    222	=> x"E4B4A696",	--mhpmcounterH7
    223	=> x"F8849E7C",	--mhpmcounterH8
    224	=> x"085E57FD",	--mhpmcounterH9
    225	=> x"076499D1",	--mhpmcounterH10
    226	=> x"A5D6B50C",	--mhpmcounterH11
    227	=> x"AE6B9B3E",	--mhpmcounterH12
    228	=> x"CCD0D516",	--mhpmcounterH13
    229	=> x"265D0119",	--mhpmcounterH14
    230	=> x"AE6ED18B",	--mhpmcounterH15
    231	=> x"C30B8E07",	--mhpmcounterH16
    232	=> x"44D80E4E",	--mhpmcounterH17
    233	=> x"8C4B52B7",	--mhpmcounterH18
    234	=> x"59A7F809",	--mhpmcounterH19
    235	=> x"11AB47E0",	--mhpmcounterH20
    236	=> x"3E6A2D93",	--mhpmcounterH21
    237	=> x"E2BB027C",	--mhpmcounterH22
    238	=> x"2E7AB1EA",	--mhpmcounterH23
    239	=> x"4C6D213A",	--mhpmcounterH24
    240	=> x"86301807",	--mhpmcounterH25
    241	=> x"9BD1C6C1",	--mhpmcounterH26
    242	=> x"247ED1D4",	--mhpmcounterH27
    243	=> x"6BFD208B",	--mhpmcounterH28
    244	=> x"FA9559C5",	--mhpmcounterH29
    245	=> x"E700B40F",	--mhpmcounterH30
    246	=> x"923C847D",	--mhpmcounterH31
    247	=> x"EDA067F5",	--mvendorid
    248	=> x"2B23F7D1",	--marchid
    249	=> x"6FB4CED8",	--mimpid
    250	=> x"76F508B6",	--mhartid
    251	=> x"05E95342",	--faulty address
    252	=> x"BC0438AF",	--faulty address
    253	=> x"604368B0",	--faulty address
    254	=> x"C122FD29",	--faulty address
    255	=> x"9BF3C712"	--faulty address
    );

--control_stim(13) = CSR_write, control_stim(12) = CSR_read, control_stim(11 downto 0) = CSR_address
constant stimulus_control : control_stim(255 downto 0) :=
    (
    0 => "1" & "0" &  x"320",	--mcountinhibit
    1 => "1" & "0" &  x"B00",	--mcycle
    2 => "1" & "0" &  x"B80",	--mcycleH
    3 => "1" & "0" &  x"B02",	--minstret
    4 => "1" & "0" &  x"B82",	--minstretH
    5 => "1" & "0" &  x"320",	--mcountinhibit
    6 => "1" & "0" &  x"300",	--mstatus
    7 => "1" & "0" &  x"304",	--mie
    8 => "1" & "0" &  x"344",	--mip
    9 => "1" & "0" &  x"305",	--mtvec
    10 => "1" & "0" &  x"340",	--mscratch
    11 => "1" & "0" &  x"341",	--mepc
    12 => "1" & "0" &  x"342",	--mcause
    13 => "1" & "0" &  x"343",	--mtval
    14 => "1" & "0" &  x"3A0",	--pmpcfg0
    15 => "1" & "0" &  x"3A1",	--pmpcfg1
    16 => "1" & "0" &  x"3A2",	--pmpcfg2
    17 => "1" & "0" &  x"3A3",	--pmpcfg3
    18 => "1" & "0" &  x"3B0",	--pmpaddr0
    19 => "1" & "0" &  x"3B1",	--pmpaddr1
    20 => "1" & "0" &  x"3B2",	--pmpaddr2
    21 => "1" & "0" &  x"3B3",	--pmpaddr3
    22 => "1" & "0" &  x"3B4",	--pmpaddr4
    23 => "1" & "0" &  x"3B5",	--pmpaddr5
    24 => "1" & "0" &  x"3B6",	--pmpaddr6
    25 => "1" & "0" &  x"3B7",	--pmpaddr7
    26 => "1" & "0" &  x"3B8",	--pmpaddr8
    27 => "1" & "0" &  x"3B9",	--pmpaddr9
    28 => "1" & "0" &  x"3BA",	--pmpaddr10
    29 => "1" & "0" &  x"3BB",	--pmpaddr11
    30 => "1" & "0" &  x"3BC",	--pmpaddr12
    31 => "1" & "0" &  x"3BD",	--pmpaddr13
    32 => "1" & "0" &  x"3BE",	--pmpaddr14
    33 => "1" & "0" &  x"3BF",	--pmpaddr15
    34	=> "1" & "0" &  x"301",	--misa
    35	=> "1" & "0" &  x"323",	--mhpmevent3
    36	=> "1" & "0" &  x"324",	--mhpmevent4
    37	=> "1" & "0" &  x"325",	--mhpmevent5
    38	=> "1" & "0" &  x"326",	--mhpmevent6
    39	=> "1" & "0" &  x"327",	--mhpmevent7
    40	=> "1" & "0" &  x"328",	--mhpmevent8
    41	=> "1" & "0" &  x"329",	--mhpmevent9
    42	=> "1" & "0" &  x"32A",	--mhpmevent10
    43	=> "1" & "0" &  x"32B",	--mhpmevent11
    44	=> "1" & "0" &  x"32C",	--mhpmevent12
    45	=> "1" & "0" &  x"32D",	--mhpmevent13
    46	=> "1" & "0" &  x"32E",	--mhpmevent14
    47	=> "1" & "0" &  x"32F",	--mhpmevent15
    48	=> "1" & "0" &  x"330",	--mhpmevent16
    49	=> "1" & "0" &  x"331",	--mhpmevent17
    50	=> "1" & "0" &  x"332",	--mhpmevent18
    51	=> "1" & "0" &  x"333",	--mhpmevent19
    52	=> "1" & "0" &  x"334",	--mhpmevent20
    53	=> "1" & "0" &  x"335",	--mhpmevent21
    54	=> "1" & "0" &  x"336",	--mhpmevent22
    55	=> "1" & "0" &  x"337",	--mhpmevent23
    56	=> "1" & "0" &  x"338",	--mhpmevent24
    57	=> "1" & "0" &  x"339",	--mhpmevent25
    58	=> "1" & "0" &  x"33A",	--mhpmevent26
    59	=> "1" & "0" &  x"33B",	--mhpmevent27
    60	=> "1" & "0" &  x"33C",	--mhpmevent28
    61	=> "1" & "0" &  x"33D",	--mhpmevent29
    62	=> "1" & "0" &  x"33E",	--mhpmevent30
    63	=> "1" & "0" &  x"33F",	--mhpmevent31
    64	=> "1" & "0" &  x"B03",	--mhpmcounter3
    65	=> "1" & "0" &  x"B04",	--mhpmcounter4
    66	=> "1" & "0" &  x"B05",	--mhpmcounter5
    67	=> "1" & "0" &  x"B06",	--mhpmcounter6
    68	=> "1" & "0" &  x"B07",	--mhpmcounter7
    69	=> "1" & "0" &  x"B08",	--mhpmcounter8
    70	=> "1" & "0" &  x"B09",	--mhpmcounter9
    71	=> "1" & "0" &  x"B0A",	--mhpmcounter10
    72	=> "1" & "0" &  x"B0B",	--mhpmcounter11
    73	=> "1" & "0" &  x"B0C",	--mhpmcounter12
    74	=> "1" & "0" &  x"B0D",	--mhpmcounter13
    75	=> "1" & "0" &  x"B0E",	--mhpmcounter14
    76	=> "1" & "0" &  x"B0F",	--mhpmcounter15
    77	=> "1" & "0" &  x"B10",	--mhpmcounter16
    78	=> "1" & "0" &  x"B11",	--mhpmcounter17
    79	=> "1" & "0" &  x"B12",	--mhpmcounter18
    80	=> "1" & "0" &  x"B13",	--mhpmcounter19
    81	=> "1" & "0" &  x"B14",	--mhpmcounter20
    82	=> "1" & "0" &  x"B15",	--mhpmcounter21
    83	=> "1" & "0" &  x"B16",	--mhpmcounter22
    84	=> "1" & "0" &  x"B17",	--mhpmcounter23
    85	=> "1" & "0" &  x"B18",	--mhpmcounter24
    86	=> "1" & "0" &  x"B19",	--mhpmcounter25
    87	=> "1" & "0" &  x"B1A",	--mhpmcounter26
    88	=> "1" & "0" &  x"B1B",	--mhpmcounter27
    89	=> "1" & "0" &  x"B1C",	--mhpmcounter28
    90	=> "1" & "0" &  x"B1D",	--mhpmcounter29
    91	=> "1" & "0" &  x"B1E",	--mhpmcounter30
    92	=> "1" & "0" &  x"B1F",	--mhpmcounter31
    93	=> "1" & "0" &  x"B83",	--mhpmcounterH3
    94	=> "1" & "0" &  x"B84",	--mhpmcounterH4
    95	=> "1" & "0" &  x"B85",	--mhpmcounterH5
    96	=> "1" & "0" &  x"B86",	--mhpmcounterH6
    97	=> "1" & "0" &  x"B87",	--mhpmcounterH7
    98	=> "1" & "0" &  x"B88",	--mhpmcounterH8
    99	=> "1" & "0" &  x"B89",	--mhpmcounterH9
    100	=> "1" & "0" &  x"B8A",	--mhpmcounterH10
    101	=> "1" & "0" &  x"B8B",	--mhpmcounterH11
    102	=> "1" & "0" &  x"B8C",	--mhpmcounterH12
    103	=> "1" & "0" &  x"B8D",	--mhpmcounterH13
    104	=> "1" & "0" &  x"B8E",	--mhpmcounterH14
    105	=> "1" & "0" &  x"B8F",	--mhpmcounterH15
    106	=> "1" & "0" &  x"B90",	--mhpmcounterH16
    107	=> "1" & "0" &  x"B91",	--mhpmcounterH17
    108	=> "1" & "0" &  x"B92",	--mhpmcounterH18
    109	=> "1" & "0" &  x"B93",	--mhpmcounterH19
    110	=> "1" & "0" &  x"B94",	--mhpmcounterH20
    111	=> "1" & "0" &  x"B95",	--mhpmcounterH21
    112	=> "1" & "0" &  x"B96",	--mhpmcounterH22
    113	=> "1" & "0" &  x"B97",	--mhpmcounterH23
    114	=> "1" & "0" &  x"B98",	--mhpmcounterH24
    115	=> "1" & "0" &  x"B99",	--mhpmcounterH25
    116	=> "1" & "0" &  x"B9A",	--mhpmcounterH26
    117	=> "1" & "0" &  x"B9B",	--mhpmcounterH27
    118	=> "1" & "0" &  x"B9C",	--mhpmcounterH28
    119	=> "1" & "0" &  x"B9D",	--mhpmcounterH29
    120	=> "1" & "0" &  x"B9E",	--mhpmcounterH30
    121	=> "1" & "0" &  x"B9F",	--mhpmcounterH31
    122	=> "1" & "0" &  x"F11",	--mvendorid
    123	=> "1" & "0" &  x"F12",	--marchid
    124	=> "1" & "0" &  x"F13",	--mimpid
    125	=> "1" & "0" &  x"F14",	--mhartid
    126	=> "0" & "1" &  x"300",	--mstatus
    127	=> "0" & "1" &  x"B82",	--minstretH
    128	=> "0" & "1" &  x"304",	--mie
    129	=> "0" & "1" &  x"305",	--mtvec
    130	=> "0" & "1" &  x"320",	--mcountinhibit
    131	=> "0" & "1" &  x"340",	--mscratch
    132	=> "0" & "1" &  x"341",	--mepc
    133	=> "0" & "1" &  x"342",	--mcause
    134	=> "0" & "1" &  x"343",	--mtval
    135	=> "0" & "1" &  x"344",	--mip
    136	=> "0" & "1" &  x"3A0",	--pmpcfg0
    137	=> "0" & "1" &  x"3A1",	--pmpcfg1
    138	=> "0" & "1" &  x"3A2",	--pmpcfg2
    139	=> "0" & "1" &  x"3A3",	--pmpcfg3
    140	=> "0" & "1" &  x"3B0",	--pmpaddr0
    141	=> "0" & "1" &  x"3B1",	--pmpaddr1
    142	=> "0" & "1" &  x"3B2",	--pmpaddr2
    143	=> "0" & "1" &  x"3B3",	--pmpaddr3
    144	=> "0" & "1" &  x"3B4",	--pmpaddr4
    145	=> "0" & "1" &  x"3B5",	--pmpaddr5
    146	=> "0" & "1" &  x"3B6",	--pmpaddr6
    147	=> "0" & "1" &  x"3B7",	--pmpaddr7
    148	=> "0" & "1" &  x"3B8",	--pmpaddr8
    149	=> "0" & "1" &  x"3B9",	--pmpaddr9
    150	=> "0" & "1" &  x"3BA",	--pmpaddr10
    151	=> "0" & "1" &  x"3BB",	--pmpaddr11
    152	=> "0" & "1" &  x"3BC",	--pmpaddr12
    153	=> "0" & "1" &  x"3BD",	--pmpaddr13
    154	=> "0" & "1" &  x"3BE",	--pmpaddr14
    155	=> "0" & "1" &  x"3BF",	--pmpaddr15
    156	=> "0" & "1" &  x"B00",	--mcycle
    157	=> "0" & "1" &  x"B02",	--minstret
    158	=> "0" & "1" &  x"B80",	--mcycleH
    159	=> "0" & "1" &  x"301",	--misa
    160	=> "0" & "1" &  x"323",	--mhpmevent3
    161	=> "0" & "1" &  x"324",	--mhpmevent4
    162	=> "0" & "1" &  x"325",	--mhpmevent5
    163	=> "0" & "1" &  x"326",	--mhpmevent6
    164	=> "0" & "1" &  x"327",	--mhpmevent7
    165	=> "0" & "1" &  x"328",	--mhpmevent8
    166	=> "0" & "1" &  x"329",	--mhpmevent9
    167	=> "0" & "1" &  x"32A",	--mhpmevent10
    168	=> "0" & "1" &  x"32B",	--mhpmevent11
    169	=> "0" & "1" &  x"32C",	--mhpmevent12
    170	=> "0" & "1" &  x"32D",	--mhpmevent13
    171	=> "0" & "1" &  x"32E",	--mhpmevent14
    172	=> "0" & "1" &  x"32F",	--mhpmevent15
    173	=> "0" & "1" &  x"330",	--mhpmevent16
    174	=> "0" & "1" &  x"331",	--mhpmevent17
    175	=> "0" & "1" &  x"332",	--mhpmevent18
    176	=> "0" & "1" &  x"333",	--mhpmevent19
    177	=> "0" & "1" &  x"334",	--mhpmevent20
    178	=> "0" & "1" &  x"335",	--mhpmevent21
    179	=> "0" & "1" &  x"336",	--mhpmevent22
    180	=> "0" & "1" &  x"337",	--mhpmevent23
    181	=> "0" & "1" &  x"338",	--mhpmevent24
    182	=> "0" & "1" &  x"339",	--mhpmevent25
    183	=> "0" & "1" &  x"33A",	--mhpmevent26
    184	=> "0" & "1" &  x"33B",	--mhpmevent27
    185	=> "0" & "1" &  x"33C",	--mhpmevent28
    186	=> "0" & "1" &  x"33D",	--mhpmevent29
    187	=> "0" & "1" &  x"33E",	--mhpmevent30
    188	=> "0" & "1" &  x"33F",	--mhpmevent31
    189	=> "0" & "1" &  x"B03",	--mhpmcounter3
    190	=> "0" & "1" &  x"B04",	--mhpmcounter4
    191	=> "0" & "1" &  x"B05",	--mhpmcounter5
    192	=> "0" & "1" &  x"B06",	--mhpmcounter6
    193	=> "0" & "1" &  x"B07",	--mhpmcounter7
    194	=> "0" & "1" &  x"B08",	--mhpmcounter8
    195	=> "0" & "1" &  x"B09",	--mhpmcounter9
    196	=> "0" & "1" &  x"B0A",	--mhpmcounter10
    197	=> "0" & "1" &  x"B0B",	--mhpmcounter11
    198	=> "0" & "1" &  x"B0C",	--mhpmcounter12
    199	=> "0" & "1" &  x"B0D",	--mhpmcounter13
    200	=> "0" & "1" &  x"B0E",	--mhpmcounter14
    201	=> "0" & "1" &  x"B0F",	--mhpmcounter15
    202	=> "0" & "1" &  x"B10",	--mhpmcounter16
    203	=> "0" & "1" &  x"B11",	--mhpmcounter17
    204	=> "0" & "1" &  x"B12",	--mhpmcounter18
    205	=> "0" & "1" &  x"B13",	--mhpmcounter19
    206	=> "0" & "1" &  x"B14",	--mhpmcounter20
    207	=> "0" & "1" &  x"B15",	--mhpmcounter21
    208	=> "0" & "1" &  x"B16",	--mhpmcounter22
    209	=> "0" & "1" &  x"B17",	--mhpmcounter23
    210	=> "0" & "1" &  x"B18",	--mhpmcounter24
    211	=> "0" & "1" &  x"B19",	--mhpmcounter25
    212	=> "0" & "1" &  x"B1A",	--mhpmcounter26
    213	=> "0" & "1" &  x"B1B",	--mhpmcounter27
    214	=> "0" & "1" &  x"B1C",	--mhpmcounter28
    215	=> "0" & "1" &  x"B1D",	--mhpmcounter29
    216	=> "0" & "1" &  x"B1E",	--mhpmcounter30
    217	=> "0" & "1" &  x"B1F",	--mhpmcounter31
    218	=> "0" & "1" &  x"B83",	--mhpmcounterH3
    219	=> "0" & "1" &  x"B84",	--mhpmcounterH4
    220	=> "0" & "1" &  x"B85",	--mhpmcounterH5
    221	=> "0" & "1" &  x"B86",	--mhpmcounterH6
    222	=> "0" & "1" &  x"B87",	--mhpmcounterH7
    223	=> "0" & "1" &  x"B88",	--mhpmcounterH8
    224	=> "0" & "1" &  x"B89",	--mhpmcounterH9
    225	=> "0" & "1" &  x"B8A",	--mhpmcounterH10
    226	=> "0" & "1" &  x"B8B",	--mhpmcounterH11
    227	=> "0" & "1" &  x"B8C",	--mhpmcounterH12
    228	=> "0" & "1" &  x"B8D",	--mhpmcounterH13
    229	=> "0" & "1" &  x"B8E",	--mhpmcounterH14
    230	=> "0" & "1" &  x"B8F",	--mhpmcounterH15
    231	=> "0" & "1" &  x"B90",	--mhpmcounterH16
    232	=> "0" & "1" &  x"B91",	--mhpmcounterH17
    233	=> "0" & "1" &  x"B92",	--mhpmcounterH18
    234	=> "0" & "1" &  x"B93",	--mhpmcounterH19
    235	=> "0" & "1" &  x"B94",	--mhpmcounterH20
    236	=> "0" & "1" &  x"B95",	--mhpmcounterH21
    237	=> "0" & "1" &  x"B96",	--mhpmcounterH22
    238	=> "0" & "1" &  x"B97",	--mhpmcounterH23
    239	=> "0" & "1" &  x"B98",	--mhpmcounterH24
    240	=> "0" & "1" &  x"B99",	--mhpmcounterH25
    241	=> "0" & "1" &  x"B9A",	--mhpmcounterH26
    242	=> "0" & "1" &  x"B9B",	--mhpmcounterH27
    243	=> "0" & "1" &  x"B9C",	--mhpmcounterH28
    244	=> "0" & "1" &  x"B9D",	--mhpmcounterH29
    245	=> "0" & "1" &  x"B9E",	--mhpmcounterH30
    246	=> "0" & "1" &  x"B9F",	--mhpmcounterH31
    247	=> "0" & "1" &  x"F11",	--mvendorid
    248	=> "0" & "1" &  x"F12",	--marchid
    249	=> "0" & "1" &  x"F13",	--mimpid
    250	=> "0" & "1" &  x"F14",	--mhartid
    251	=> "1" & "1" &  x"FFF",	--faulty address
    252	=> "1" & "0" &  x"DEA",	--faulty address
    253	=> "1" & "0" &  x"754",	--faulty address
    254	=> "0" & "1" &  x"193",	--faulty address
    255	=> "0" & "0" &  x"C23"	--faulty address
    );
end package;
